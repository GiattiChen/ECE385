module wall(input [9:0] wallX,
				input [9:0] wallY,
				input [7:0] p1ab,
				input logic isDoor,
				output logic [2:0] cidx
				);
			
	
	logic [2:0] IMG [899:0] = '{3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b010,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b001,3'b000,3'b000,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b010,3'b010,3'b010,3'b010,3'b010,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b010,3'b000,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b001,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b010,3'b001,3'b010,3'b000,3'b010,3'b010,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b000,3'b000,3'b001,3'b010,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b010,3'b001,3'b010,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b001,3'b010,3'b001,3'b010,3'b001,3'b001,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b010,3'b010,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b000,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b010,3'b000,3'b001,3'b000,3'b000,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b010,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b010,3'b010,3'b000,3'b000,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b000,3'b000,3'b000,3'b000,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b000,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b001,3'b000,3'b001,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b001,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b000,3'b000,3'b010,3'b000,3'b000,3'b001,3'b001,3'b010,3'b000,3'b001,3'b001,3'b001,3'b010,3'b000,3'b010,3'b010,3'b000,3'b001,3'b001,3'b000,3'b001,3'b001,3'b010};	
	logic	DOOR[899:0] = '{0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic [9:0] idx;
	assign idx = wallX*30 + wallY;
	always_comb
		begin
			if (p1ab == 1 && isDoor == 1 && DOOR[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else
				begin
					cidx = IMG[899 - idx];
				end
		end
endmodule


module road(input [9:0] roadX,
				input [9:0] roadY,
				input [7:0] p1ab,
				input [7:0] p2ab,
				input [1:0] SD,
				output logic [2:0] cidx
				);
			
	
	logic [2:0] IMG1 [899:0] = '{3'b100,3'b101,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b101,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b101,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b101,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b101,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b101,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b101,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b101,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b101,3'b101,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b101,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b101,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b101,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b101,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b110,3'b100,3'b110,3'b101,3'b110,3'b100,3'b100,3'b110,3'b110,3'b110,3'b110,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b101,3'b100,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b110,3'b110,3'b100,3'b100,3'b100,3'b100,3'b100,3'b110,3'b100,3'b110,3'b100};	
	logic SHIT[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic PLANES[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic PLANED[899:0] = '{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	logic [9:0] idx;
	assign idx = roadX*30 + roadY;
		always_comb
		begin
			cidx = IMG1[899 - idx];
			if (p1ab == 0 && SD == 2 && PLANES[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else if (p1ab == 0 && SD == 3 && PLANED[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
			else if (p2ab == 1 && SD == 1 && SHIT[899 -idx] == 1)
				begin
					cidx = 3'b111;
				end
		end
endmodule

module big(input [9:0] nX,
				input [9:0] nY,
				output logic [10:0] cidx
				);
	logic [9:0] IMG [24999:0] = '{155,83,147,155,228,155,155,227,293,221,220,220,156,292,220,220,220,229,156,156,220,156,155,155,292,220,220,156,291,156,219,293,355,427,427,355,363,428,419,355,419,419,354,355,419,419,419,419,419,419,354,419,355,354,354,291,419,419,355,355,355,155,147,219,355,147,355,419,355,419,146,74,419,290,419,355,211,427,354,354,419,418,419,355,354,346,419,282,282,146,354,354,211,73,0,136,144,65,74,209,73,145,1,0,72,0,72,81,74,0,73,73,137,72,145,64,0,73,137,137,136,73,137,1,64,228,155,82,147,82,293,155,154,155,292,220,292,155,220,219,220,292,292,220,156,156,155,156,156,156,356,156,220,156,228,220,302,229,219,147,364,356,292,292,219,74,147,74,147,156,147,147,147,146,147,147,138,147,219,146,148,74,147,147,147,147,83,147,147,147,83,147,219,74,291,147,2,282,290,354,145,147,354,354,419,283,210,419,147,355,419,283,219,155,73,219,346,74,1,0,73,137,1,137,73,1,64,1,65,73,0,0,73,73,1,73,73,73,72,144,64,73,73,137,73,137,65,73,0,0,156,229,219,155,83,147,156,155,155,155,228,356,228,220,292,220,292,229,228,147,220,220,155,155,155,147,356,220,294,294,292,220,293,156,229,219,292,221,220,356,365,147,147,147,147,83,156,147,219,219,148,146,83,147,74,83,84,292,147,156,156,147,83,147,74,74,155,148,146,155,74,1,290,362,354,146,283,290,427,355,156,219,355,283,282,419,291,74,146,219,147,219,65,1,0,1,73,1,73,73,1,64,65,73,73,0,73,72,0,1,73,73,138,64,136,73,65,73,64,1,145,65,73,65,64,219,219,221,156,219,155,155,209,218,155,228,228,155,301,292,220,220,220,229,148,220,293,219,155,163,294,227,227,156,293,302,292,364,147,221,156,364,229,220,293,155,73,147,147,147,82,84,83,147,220,220,147,146,148,147,83,148,148,155,148,148,156,147,147,147,137,148,82,219,73,10,65,281,362,290,291,147,362,419,283,155,219,218,147,219,219,83,156,147,147,73,219,283,1,65,1,73,1,137,65,1,73,65,73,73,0,0,72,0,1,64,145,73,145,64,64,65,73,64,73,73,65,73,66,1,147,156,220,220,156,75,74,155,137,282,282,155,228,220,220,365,220,364,221,229,220,221,302,292,156,155,228,163,227,156,220,356,292,292,147,220,355,219,221,211,283,74,83,147,74,147,147,220,211,147,147,292,147,220,156,82,84,156,147,148,157,83,74,147,82,146,83,155,219,146,10,281,362,291,355,355,219,355,419,220,219,155,155,147,292,219,147,83,83,147,283,147,219,74,65,65,65,73,73,1,1,73,1,73,73,0,64,137,1,0,73,144,145,136,72,145,65,0,65,137,74,137,73,137,1,75,75,83,148,155,227,75,76,219,210,210,282,219,156,220,220,365,229,293,293,220,220,293,219,156,156,292,227,155,220,219,292,292,292,293,292,218,355,156,220,147,220,84,147,147,156,293,292,147,364,364,363,363,148,292,147,83,147,219,83,1,156,147,147,9,73,65,155,220,74,83,137,428,354,292,355,155,428,419,147,219,147,156,219,83,155,82,83,75,147,219,83,219,74,66,65,1,73,73,73,73,73,73,73,73,0,73,73,73,65,73,136,73,137,137,137,73,64,137,137,65,138,65,137,1,75,75,75,74,75,147,156,155,76,148,219,209,282,282,220,156,220,365,229,364,364,220,148,228,147,157,220,146,227,156,228,228,292,356,211,364,301,356,292,365,293,221,83,147,220,147,301,211,364,502,438,365,291,364,228,147,155,147,219,221,73,148,74,156,147,82,146,83,220,147,355,74,227,355,155,364,147,291,355,156,219,74,220,355,147,155,147,75,74,147,83,219,219,74,1,65,1,1,73,9,73,73,1,73,0,73,65,8,1,0,147,137,74,145,145,64,137,73,137,74,137,137,1,1,1,211,83,11,75,75,75,75,156,156,291,302,221,210,274,293,293,292,221,229,293,292,220,220,75,147,147,156,291,292,228,221,292,221,293,365,292,220,301,355,293,293,228,155,156,156,220,219,438,364,365,437,429,365,355,430,147,220,84,155,220,1,156,83,148,156,75,155,148,156,147,291,290,291,292,220,355,155,156,219,148,220,219,220,283,155,155,82,83,82,75,74,283,218,220,74,1,0,73,73,65,1,73,73,1,65,9,65,145,73,0,210,137,74,145,145,137,65,137,136,74,74,201,73,1,137,146,147,147,75,83,147,147,147,83,147,220,302,294,291,210,283,366,220,156,229,365,365,221,147,147,220,146,220,292,283,220,220,229,221,366,292,229,365,292,364,365,229,156,220,148,292,156,427,437,365,291,373,437,364,155,218,148,148,220,147,229,148,83,155,220,148,220,83,220,75,355,427,227,292,156,291,219,148,219,220,292,219,292,292,219,83,147,83,147,74,147,220,292,147,282,65,73,0,73,73,72,73,73,1,0,73,1,74,73,0,145,144,145,137,145,137,0,137,64,73,74,137,65,138,1,147,147,156,84,147,84,148,147,219,75,156,228,293,302,283,209,365,292,219,156,221,293,293,221,220,147,148,292,220,364,220,155,228,147,293,365,221,229,366,364,365,229,228,147,148,220,293,364,373,510,364,291,501,220,219,74,157,229,156,84,148,147,156,220,228,83,284,147,292,147,291,355,283,292,156,355,146,147,219,147,220,283,147,291,292,83,219,83,147,83,10,83,292,83,283,73,75,73,65,73,73,137,73,73,0,1,1,74,0,0,144,72,137,74,73,73,137,137,73,137,73,137,137,137,73,83,75,84,147,76,83,147,84,84,212,147,155,221,293,221,292,283,282,282,218,282,292,365,302,229,83,148,82,220,293,292,292,228,293,293,292,364,156,366,292,365,294,365,220,156,148,220,220,365,438,438,227,355,228,366,147,84,220,1,156,84,75,82,156,219,83,220,227,228,146,363,363,220,292,220,356,146,229,219,219,291,219,283,356,227,147,147,147,155,147,75,74,292,148,291,74,75,10,0,72,73,1,73,1,9,73,2,75,74,0,144,74,145,146,74,137,137,73,74,137,65,73,138,137,138,83,83,83,84,83,84,147,84,148,83,147,84,75,156,148,229,221,283,274,292,210,429,365,374,293,220,84,83,74,292,364,229,220,229,293,366,357,228,293,430,292,229,291,292,228,220,219,438,220,293,228,156,147,220,147,155,148,83,74,156,148,156,83,83,146,148,211,227,228,292,363,355,356,292,292,356,364,220,228,219,219,219,228,155,228,219,147,146,219,146,83,147,220,147,219,75,74,75,1,65,73,1,74,65,73,73,65,75,73,1,72,146,144,73,74,137,137,1,73,137,1,137,0,0,1,84,147,148,147,148,148,147,148,156,84,219,148,83,147,149,220,228,293,283,218,357,428,229,365,429,229,156,84,83,227,229,356,220,229,221,219,439,228,365,366,219,293,293,219,155,155,219,219,228,147,210,365,293,155,211,156,156,147,156,156,156,74,74,147,219,138,284,291,220,220,364,291,363,356,227,356,364,228,228,364,220,219,219,219,155,220,155,292,292,219,147,219,155,147,155,75,147,75,74,66,74,1,146,9,72,9,1,65,75,65,0,145,144,64,65,65,65,1,73,137,137,0,0,64,1,84,76,83,147,75,84,83,83,148,147,147,147,74,75,156,76,228,302,301,210,284,282,220,229,356,429,284,147,148,83,229,229,365,220,229,220,366,229,356,292,366,147,293,430,228,284,156,219,220,83,156,219,156,156,147,156,156,220,156,83,156,229,74,83,147,146,147,291,228,156,427,219,362,354,291,291,355,364,291,364,292,292,156,292,147,355,219,292,219,228,219,355,228,147,147,147,74,75,75,73,74,65,0,9,73,73,1,0,74,0,64,74,81,64,73,145,2,0,0,0,72,0,64,0,0,84,76,148,83,147,83,220,84,147,156,148,147,74,73,74,220,148,293,293,301,209,301,282,228,365,356,293,292,157,147,74,229,300,228,228,228,219,365,229,356,366,292,293,438,356,147,83,75,147,75,148,73,155,83,147,148,220,228,156,221,156,220,74,73,156,147,146,291,219,147,428,291,291,363,363,291,292,364,364,364,365,292,220,220,219,219,292,292,220,292,228,292,83,219,156,211,75,76,82,74,65,74,0,81,73,73,73,0,1,1,137,1,137,146,66,1,74,138,146,145,2,72,72,136,1,84,148,84,148,147,211,75,147,147,148,147,147,148,73,9,146,220,302,293,302,228,274,273,283,229,356,293,220,293,221,74,74,292,293,228,293,365,364,229,228,364,292,293,366,363,219,220,156,74,148,83,148,156,147,156,147,148,147,156,156,221,220,148,73,156,148,74,210,291,147,356,291,228,363,363,362,363,428,364,364,292,155,292,155,219,156,356,292,292,83,292,219,75,220,156,211,75,147,74,0,1,1,73,73,2,65,0,0,0,73,210,1,74,65,1,2,2,73,210,137,65,72,136,0,144,148,220,84,84,147,147,155,148,148,148,156,74,156,74,73,73,219,220,291,365,229,283,282,283,293,302,293,365,221,229,74,74,291,302,293,293,292,356,229,229,291,230,293,221,291,219,74,221,138,220,220,157,156,220,156,292,148,155,220,156,221,156,148,147,156,156,220,220,147,73,219,219,300,228,363,371,363,300,364,364,365,156,364,292,155,220,220,364,292,83,228,219,83,220,156,291,82,74,74,65,74,0,9,73,75,73,73,73,72,137,217,73,138,73,1,74,74,73,137,210,1,65,144,0,144,157,83,148,148,76,147,147,76,148,75,156,221,84,146,149,137,82,292,283,283,292,220,282,302,283,229,366,221,292,229,229,74,155,294,230,229,293,292,292,228,292,294,292,293,283,156,82,147,220,147,147,148,148,228,220,219,156,220,156,157,221,220,157,219,156,147,283,220,83,74,83,283,219,292,228,364,363,363,364,364,292,364,155,291,292,156,74,228,364,210,75,220,83,155,291,210,75,75,75,74,1,0,1,0,1,0,72,73,64,64,145,73,137,73,146,138,74,73,137,210,65,64,144,1,136,84,84,147,148,148,84,147,74,219,156,148,156,220,84,73,221,219,138,220,282,428,294,366,302,210,293,293,221,293,229,221,74,146,356,229,228,221,293,293,365,364,294,293,293,219,220,219,156,147,156,157,148,156,219,156,220,220,155,155,156,221,219,156,147,148,83,147,156,75,74,74,219,147,365,228,220,364,363,292,292,291,364,364,220,291,155,147,147,292,364,147,83,148,220,364,138,75,211,75,146,0,73,9,72,64,73,145,1,73,64,145,73,146,74,146,138,2,137,73,146,146,65,72,1,73,84,84,84,147,148,75,148,229,148,220,75,74,155,147,210,148,74,75,220,292,292,366,366,283,302,283,293,301,294,229,221,75,74,292,293,292,156,228,293,293,364,294,293,293,292,155,147,148,74,147,156,156,156,155,155,220,228,155,147,83,229,155,156,148,83,156,83,156,10,83,83,11,83,228,365,228,301,365,363,292,428,291,292,292,220,291,155,146,147,292,147,74,83,292,364,147,74,75,147,73,1,0,8,73,0,73,74,1,74,145,136,137,137,138,74,146,10,73,137,145,218,0,136,73,136,148,149,75,83,147,147,84,227,76,283,147,82,147,220,220,73,147,147,82,220,229,365,367,284,221,282,293,229,293,293,221,156,219,292,293,357,229,220,357,293,365,229,364,294,294,220,147,155,147,156,283,362,209,363,427,289,146,290,219,146,156,292,156,83,147,84,156,147,221,83,148,75,83,220,364,301,292,292,218,363,363,364,355,365,228,220,300,291,74,156,292,83,147,156,292,75,74,75,74,0,1,1,145,73,0,74,74,73,73,75,74,2,65,74,73,74,74,73,137,146,145,137,0,0,0,156,84,147,84,156,283,83,155,84,147,220,220,74,147,149,73,138,147,148,283,229,367,366,293,284,283,292,294,293,220,148,148,219,219,293,293,156,221,366,293,294,230,363,229,294,291,83,220,156,220,209,363,363,290,291,236,363,362,354,146,219,156,228,148,156,156,156,147,148,83,10,84,75,220,156,292,291,300,356,292,363,292,428,300,292,220,220,156,291,83,228,300,147,156,220,75,139,74,74,0,73,1,145,73,73,74,10,211,74,74,74,74,73,137,74,146,138,146,146,137,210,209,73,0,72,147,148,148,84,74,220,148,147,74,147,147,148,220,147,148,146,74,73,149,293,292,367,294,292,210,284,292,284,356,211,148,148,154,220,293,220,292,293,366,229,302,302,364,293,220,291,156,220,156,147,290,299,363,363,372,363,436,299,363,354,354,156,156,148,148,92,83,148,220,220,74,156,75,148,148,156,228,364,292,356,364,292,291,292,292,292,220,156,228,147,155,364,83,83,292,74,74,75,73,1,65,1,73,73,76,73,10,73,73,73,74,73,146,210,82,73,74,73,137,210,145,282,0,136,136,148,148,149,83,82,74,147,148,156,147,147,147,156,83,148,84,147,73,148,292,291,302,229,364,209,220,220,220,220,220,148,148,299,292,293,293,365,365,302,293,293,294,364,220,293,219,157,220,290,363,373,362,436,436,436,427,363,435,363,363,352,220,156,156,156,220,147,148,84,292,147,147,83,75,156,220,292,292,291,228,429,363,228,220,156,292,292,220,292,148,292,365,82,83,147,74,75,75,0,73,73,73,73,0,74,146,10,65,0,0,0,0,0,0,0,64,64,137,137,145,145,201,0,208,0,220,84,83,83,147,156,156,147,147,147,156,292,83,221,156,157,156,146,83,75,291,220,292,364,210,292,221,293,292,364,293,292,291,293,293,293,293,364,302,220,293,294,365,220,230,366,157,157,289,362,300,362,436,363,436,435,363,372,372,354,363,365,156,157,148,155,292,156,157,147,156,83,84,355,147,148,220,228,220,228,428,364,219,220,148,292,292,228,156,83,147,364,219,147,220,75,75,138,1,73,73,1,2,65,73,0,0,0,0,0,64,64,128,64,64,64,64,0,64,0,73,72,0,0,1,75,84,148,147,148,147,156,292,156,83,148,156,147,149,156,148,294,220,146,147,283,292,429,219,292,292,221,221,229,429,293,221,219,220,366,293,365,365,294,366,302,293,292,293,230,155,157,157,227,289,283,372,362,502,490,501,426,371,291,363,292,237,156,156,220,156,220,147,148,148,156,228,84,148,220,148,148,228,220,292,364,292,228,292,156,292,364,292,156,220,147,220,292,292,356,76,75,73,64,146,74,138,147,0,73,64,0,0,0,0,0,0,0,0,0,0,0,0,64,64,0,64,64,0,0,75,147,148,211,219,148,147,156,156,83,220,157,147,148,149,148,148,221,147,148,146,293,364,218,293,282,293,220,293,365,366,429,293,357,366,293,293,364,294,366,302,293,293,294,229,156,156,291,300,362,436,436,426,501,510,510,427,436,427,362,354,219,156,156,84,75,293,83,228,147,148,156,83,83,220,155,148,220,220,228,291,356,292,292,148,292,364,155,220,155,219,156,292,228,292,76,75,0,73,64,137,64,0,0,0,72,64,136,0,0,0,0,0,0,0,0,0,0,0,0,0,0,64,64,0,156,147,84,148,147,147,148,148,147,148,75,83,147,84,148,147,147,156,156,147,147,294,355,227,293,283,229,229,292,292,365,365,293,302,293,293,293,364,293,365,294,156,292,220,229,156,156,290,364,289,300,436,426,425,425,363,428,363,362,362,361,228,228,147,75,75,220,148,155,156,147,83,74,74,83,147,148,220,292,219,283,210,219,292,147,292,291,156,156,156,355,220,292,83,220,147,75,1,65,64,64,145,0,64,0,64,0,0,0,0,64,64,64,64,64,64,64,64,64,128,128,64,0,0,64,74,155,156,148,147,156,84,139,147,148,76,149,147,148,156,148,83,83,148,83,83,230,355,292,292,146,220,293,292,292,365,501,301,293,293,293,356,364,301,292,364,157,292,292,148,83,219,82,282,146,362,291,362,435,363,300,363,372,236,227,300,220,228,147,147,65,64,64,128,354,64,137,209,64,0,0,64,64,137,73,137,146,145,136,82,219,282,291,219,155,356,156,292,148,219,147,75,0,73,65,209,136,64,64,0,0,0,64,0,0,0,0,0,0,0,0,0,128,64,64,64,64,64,64,64,75,147,148,148,76,148,147,75,

84,148,147,148,83,147,148,147,148,156,148,157,74,229,364,364,364,210,220,156,210,137,137,137,64,73,72,72,72,64,64,73,72,146,282,137,146,73,64,65,146,353,299,364,363,363,362,362,372,362,372,299,146,129,128,128,64,0,0,0,0,0,0,0,0,0,0,0,0,64,64,64,64,64,0,72,146,137,0,73,146,155,291,156,228,219,155,147,73,137,73,137,64,0,0,0,0,0,0,0,0,0,64,64,64,64,0,0,64,0,0,0,136,64,64,64,64,147,83,148,147,148,147,156,220,148,149,83,84,83,147,220,147,147,157,156,157,147,220,293,364,292,155,220,221,293,292,220,292,283,146,137,136,64,64,0,0,72,0,0,0,64,64,72,72,8,72,64,0,145,290,363,291,283,209,128,136,128,128,128,128,128,128,0,64,64,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,64,0,0,145,73,73,73,1,1,0,65,0,64,0,0,0,0,0,0,0,64,64,64,0,64,72,0,0,0,0,0,0,64,0,72,0,0,136,219,75,148,147,75,155,156,156,148,157,75,156,147,83,148,76,74,157,156,221,83,293,302,366,293,219,220,302,228,302,229,293,293,293,229,292,292,283,136,128,136,8,8,0,0,0,0,64,136,201,137,72,73,0,0,65,73,282,428,210,200,128,128,0,8,0,128,128,64,64,64,0,0,0,0,0,0,0,0,0,0,0,0,64,0,0,0,0,0,0,0,0,64,128,64,128,64,0,0,0,0,0,0,0,72,128,128,64,0,64,64,0,0,0,0,0,0,0,0,64,0,0,64,0,0,283,76,147,148,148,155,148,156,148,157,147,220,148,83,220,76,75,148,83,157,282,367,228,302,228,220,302,302,229,302,156,229,294,302,293,292,230,292,220,291,137,136,136,72,72,0,64,128,64,0,0,0,64,72,137,72,64,0,64,64,136,64,64,273,201,136,0,0,0,64,128,128,128,64,0,0,0,0,0,0,0,0,0,0,0,0,0,64,0,0,0,0,64,0,0,0,0,0,0,0,0,0,64,136,128,128,64,64,64,64,64,64,64,64,0,0,0,0,0,0,0,0,0,0,0,211,76,83,148,156,155,148,156,148,148,75,156,157,83,155,75,74,148,83,75,283,294,220,293,220,293,293,302,357,294,220,293,294,229,294,292,293,220,220,156,219,72,72,64,0,0,0,0,0,0,0,0,64,0,64,72,64,128,200,136,0,0,64,0,0,64,128,128,128,0,0,0,0,0,0,0,0,8,0,8,0,0,0,0,0,0,0,137,0,0,0,0,145,136,128,128,128,64,64,64,64,64,64,64,209,64,0,0,8,0,0,0,0,0,64,64,128,64,0,0,0,0,0,64,0,147,147,147,147,156,219,211,148,220,84,148,156,148,156,74,147,147,83,211,147,292,229,220,302,293,302,293,365,293,293,283,293,283,292,293,292,292,293,291,200,136,137,73,74,136,136,128,128,128,128,128,128,128,128,128,128,64,64,64,0,8,0,0,0,72,0,0,64,136,200,128,64,0,0,0,0,0,0,0,0,0,0,0,0,0,73,0,0,0,0,0,0,0,0,0,72,64,0,0,0,8,0,0,210,0,0,0,0,0,0,0,0,0,0,0,0,64,64,64,64,0,0,0,209,64,211,147,211,147,146,219,219,155,147,147,284,156,147,147,83,83,148,219,147,283,220,293,156,229,229,294,229,365,201,136,210,137,136,128,136,136,128,128,136,136,73,72,72,72,72,72,72,72,72,8,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,128,128,200,128,128,128,128,64,0,0,0,0,0,0,0,0,0,0,73,0,0,0,0,0,0,72,72,72,0,0,0,0,0,0,0,0,0,0,64,136,0,0,0,0,0,0,0,0,0,0,64,0,0,0,8,64,137,137,137,136,136,136,136,64,64,72,64,72,72,64,64,72,74,146,147,355,220,229,228,228,293,229,365,366,292,73,8,73,72,145,73,72,9,9,8,8,8,9,8,73,73,73,72,8,8,8,72,8,8,8,8,8,64,64,0,64,0,0,0,0,0,0,0,0,0,0,64,128,128,128,72,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,136,136,137,0,0,64,0,0,0,72,72,73,0,0,0,0,0,0,64,64,0,0,0,0,0,0,0,0,137,64,64,72,0,0,64,64,72,64,72,72,73,64,64,72,72,72,8,73,73,73,72,72,64,72,136,210,364,292,292,364,146,209,64,64,64,64,64,64,136,128,128,128,128,128,128,64,72,64,64,64,64,64,64,64,64,0,72,8,0,72,8,0,0,72,0,8,0,0,0,0,0,0,0,0,0,0,0,201,128,128,137,64,128,128,136,137,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,64,0,0,0,0,0,72,64,0,0,0,0,0,0,0,0,0,64,64,0,0,72,8,72,72,0,72,72,72,136,137,137,137,137,136,136,136,136,72,73,72,64,72,64,64,72,137,72,64,64,64,136,64,73,8,8,72,64,64,64,64,64,0,8,8,72,72,136,128,128,128,128,128,128,64,64,64,64,64,64,64,64,64,0,0,0,0,0,64,0,64,64,0,0,64,0,64,64,128,128,128,200,64,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,72,64,0,0,0,0,0,0,145,0,0,64,0,0,72,0,0,0,0,0,0,0,0,0,0,72,0,136,137,137,137,146,147,155,220,147,148,148,156,148,83,147,74,146,137,137,72,8,72,72,136,136,72,145,72,72,8,8,9,8,8,8,9,8,72,8,64,0,8,8,8,9,8,8,8,0,64,64,64,128,200,137,64,64,64,64,64,64,64,64,128,72,0,64,0,0,64,64,64,64,64,0,0,72,64,0,0,0,0,0,0,0,0,0,0,64,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,136,72,0,218,0,0,0,0,0,0,210,0,64,64,0,0,0,0,210,211,291,281,355,291,502,437,219,301,220,147,147,157,149,157,220,147,356,218,136,136,72,72,9,9,9,8,9,8,8,8,73,145,73,218,218,8,8,9,9,9,8,8,8,8,8,8,8,8,8,64,0,0,0,0,0,8,72,0,64,64,64,64,72,8,0,0,0,0,0,0,0,0,64,137,0,0,0,0,0,0,64,0,0,0,0,0,0,0,64,64,0,0,0,0,0,0,0,0,282,0,0,0,0,0,0,64,64,145,0,0,0,0,0,0,0,0,0,0,0,0,0,137,0,357,502,218,354,437,291,363,427,354,283,301,219,83,156,84,84,157,283,221,292,364,209,136,72,72,72,8,8,0,0,0,0,0,8,8,8,9,8,9,8,8,8,0,0,0,8,8,8,8,209,72,0,0,0,0,8,0,8,0,0,8,8,0,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,0,0,0,0,72,128,128,64,64,0,0,0,0,64,128,72,0,0,64,0,0,0,0,0,64,64,209,0,0,0,281,136,64,72,73,0,72,0,0,0,64,0,64,64,0,0,0,427,355,510,355,364,437,425,427,353,362,292,219,156,148,157,156,157,364,230,221,229,356,291,209,137,73,73,81,8,64,72,72,64,64,64,64,64,0,0,0,8,145,145,72,8,72,145,73,8,8,8,8,0,0,8,0,0,72,0,0,0,72,64,72,0,0,0,0,0,9,8,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,137,72,64,64,64,64,128,128,64,209,0,0,0,0,0,0,0,136,136,128,128,128,128,200,128,128,64,128,64,64,209,128,0,64,64,0,0,0,64,219,365,283,428,425,362,361,354,353,291,426,365,157,148,157,156,158,292,157,221,302,429,293,293,292,145,210,72,64,64,0,65,64,64,64,64,136,136,273,137,136,64,137,72,72,72,0,8,0,8,72,72,72,0,0,72,73,72,8,72,0,0,0,8,0,0,8,0,72,8,8,73,8,64,0,291,0,0,0,0,0,0,0,0,0,0,0,0,0,281,200,200,128,128,64,64,136,64,128,64,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,72,64,64,64,64,0,0,0,0,0,290,363,364,427,510,428,426,437,354,362,363,502,156,148,156,220,229,302,230,302,366,291,302,430,292,301,428,428,364,293,364,292,428,292,365,356,283,292,219,283,210,146,74,73,73,73,8,8,8,8,0,0,8,0,0,0,0,0,0,0,64,64,64,64,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,0,0,0,0,137,201,136,128,128,128,128,273,64,0,0,0,0,0,0,64,64,128,136,0,0,0,0,0,354,64,0,0,0,8,72,64,64,64,64,0,0,72,0,0,0,0,363,363,436,363,498,498,425,498,362,425,427,292,157,148,147,156,293,148,220,366,292,301,366,437,229,365,293,293,293,367,292,229,293,365,366,293,366,301,220,156,229,147,219,220,155,73,82,74,74,74,73,72,0,8,8,72,136,209,64,64,0,0,0,64,64,64,64,64,64,0,72,8,72,72,137,9,0,0,0,0,0,64,128,128,128,64,64,64,64,0,128,64,0,0,0,0,0,0,0,64,64,64,0,0,0,0,0,0,0,73,8,0,64,64,64,0,0,136,0,64,0,0,64,64,0,216,363,363,425,489,497,490,490,426,436,354,219,157,220,148,221,364,84,292,366,293,229,365,366,365,156,291,302,228,367,293,229,429,366,292,366,293,229,157,229,156,147,156,83,219,128,136,128,128,136,136,128,128,128,200,128,200,136,72,64,64,64,0,0,0,0,0,0,8,0,72,8,8,0,8,8,0,0,72,128,128,64,0,0,8,0,0,0,64,64,64,72,0,64,64,0,0,0,0,0,0,64,136,136,72,0,0,0,0,64,0,0,64,64,64,0,0,64,0,64,64,354,64,0,0,363,354,364,490,489,417,489,489,353,437,354,219,157,220,82,157,220,156,365,366,156,301,438,375,293,228,220,293,220,367,293,292,366,367,293,375,293,157,147,220,157,365,155,147,155,74,64,137,64,64,64,64,64,64,64,64,64,64,128,64,64,64,64,64,136,72,136,64,72,8,0,8,8,8,8,64,273,273,136,72,72,72,0,0,0,0,0,64,8,0,0,282,136,0,0,64,0,0,0,0,0,0,273,128,64,64,64,64,0,0,64,64,64,0,0,64,0,64,64,64,0,0,0,0,0,291,290,437,490,489,425,425,489,354,363,354,292,230,149,148,157,156,229,366,366,293,430,365,302,220,356,302,283,366,302,292,429,293,302,301,375,229,156,74,156,293,292,157,429,155,156,429,147,147,74,293,220,292,292,292,428,0,73,219,155,220,220,147,73,73,137,146,137,136,72,72,72,72,72,64,72,64,0,64,136,128,128,200,128,200,128,128,136,136,209,64,0,0,72,64,64,64,0,64,0,0,0,0,64,128,136,0,136,64,64,64,64,0,0,0,0,0,0,0,0,0,8,0,0,0,283,354,501,499,497,489,489,498,429,427,437,438,221,156,156,220,229,229,293,294,156,292,366,229,283,367,365,228,437,301,292,365,229,301,366,301,157,74,147,157,301,148,148,156,1,147,83,147,74,229,156,229,156,228,293,1,147,156,156,156,157,221,148,83,156,221,156,146,156,155,283,282,346,64,0,0,0,64,0,0,64,0,64,64,64,8,8,72,0,0,0,136,64,0,0,0,0,0,0,64,64,0,0,64,128,128,128,209,136,64,64,64,64,64,72,0,136,0,0,0,64,72,0,0,0,228,436,436,363,426,434,426,361,427,363,364,439,157,156,229,365,229,374,366,293,229,293,229,228,292,375,228,374,365,292,292,294,293,374,366,294,147,155,156,301,220,156,364,147,156,292,156,74,156,146,74,147,83,365,74,0,165,228,156,229,229,157,156,229,221,228,220,82,148,156,284,220,228,356,81,82,155,146,154,145,81,8,72,72,0,0,0,0,0,0,0,64,64,64,64,64,136,0,0,136,64,0,64,0,0,128,128,128,64,64,64,0,0,0,0,0,0,0,0,128,64,0,0,0,0,355,291,428,427,354,435,373,

363,363,364,362,220,148,220,156,220,365,366,293,365,293,366,228,302,366,301,366,374,228,291,293,294,438,439,366,229,293,156,229,156,293,292,83,229,228,156,0,73,83,0,148,74,229,219,0,156,156,156,156,229,157,147,229,230,220,229,156,147,156,74,147,229,155,292,73,220,155,146,72,64,0,0,0,64,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,64,64,136,64,72,137,128,128,136,64,145,136,72,209,209,201,128,128,128,128,64,64,0,0,64,128,437,436,354,426,354,363,426,426,364,290,291,157,148,221,156,147,366,367,302,292,367,229,293,292,365,292,438,292,292,357,293,301,439,374,221,366,365,156,156,156,220,156,9,83,147,147,147,74,137,83,147,84,293,73,74,220,228,156,156,302,229,156,293,302,156,229,147,228,228,220,229,292,209,137,73,73,65,64,64,64,0,0,0,0,72,0,0,64,0,128,64,128,64,136,128,0,0,0,64,0,137,64,64,0,0,283,64,64,0,0,64,64,64,64,64,64,64,0,0,0,0,0,0,128,0,147,219,364,355,219,428,356,292,439,366,157,156,149,147,75,293,293,293,293,367,302,292,291,356,301,365,292,229,293,219,293,439,439,301,229,292,0,147,75,74,156,156,0,73,148,228,147,147,156,157,157,220,301,147,220,229,229,156,229,301,147,229,302,220,156,229,74,155,9,147,228,73,74,0,73,9,73,82,73,73,81,9,73,81,73,145,72,72,72,64,136,128,72,0,0,0,64,64,64,64,64,0,0,0,0,0,64,128,72,64,0,0,0,0,0,0,0,0,0,209,64,64,64,0,0,148,83,148,229,237,365,366,156,156,156,157,156,157,75,148,293,220,366,229,293,293,294,292,365,374,292,228,292,293,365,439,438,356,294,155,0,0,75,74,10,156,72,64,229,147,229,148,294,157,292,148,293,220,164,293,229,156,148,302,293,156,229,365,148,229,365,74,156,219,9,220,228,74,220,147,228,219,156,229,83,156,74,155,147,147,82,74,146,219,146,64,0,0,64,0,0,0,64,64,0,0,0,0,0,72,0,72,128,128,72,209,209,8,0,0,0,0,0,0,64,128,64,0,0,0,148,76,221,148,157,220,221,148,157,156,149,148,157,139,229,302,293,293,229,229,302,357,438,366,366,365,293,366,294,228,365,365,302,292,145,146,229,228,9,83,147,0,137,229,1,74,156,83,229,147,293,229,229,228,156,157,156,229,292,156,220,228,156,229,301,147,219,9,147,220,74,228,64,229,147,228,220,157,147,156,147,147,147,74,73,1,73,147,147,219,220,219,64,0,0,64,64,0,0,0,64,64,64,64,136,137,144,346,128,64,0,0,0,0,136,72,0,72,0,0,64,0,0,8,136,148,148,148,148,148,220,156,148,156,75,221,156,221,292,293,294,366,229,221,293,293,439,429,365,366,364,365,375,156,228,367,302,228,156,74,83,147,146,73,9,73,74,220,147,74,156,220,156,148,220,220,293,221,164,229,220,156,156,301,366,366,511,228,229,365,219,438,74,147,292,228,220,147,292,219,292,83,155,1,64,0,0,0,0,0,0,0,0,0,1,147,219,218,74,64,0,0,0,0,0,0,0,209,209,136,64,64,64,64,128,64,136,72,0,0,0,0,0,64,64,0,0,64,64,64,148,147,148,156,149,156,221,149,156,221,149,83,293,229,147,293,292,229,302,365,439,365,437,366,436,437,294,303,229,375,294,156,156,75,229,228,148,74,74,74,64,219,0,219,147,229,157,293,229,229,156,294,229,229,156,357,156,301,228,147,228,291,439,357,356,291,219,74,292,292,229,146,229,293,155,291,64,0,0,64,136,72,0,0,0,64,64,128,136,64,0,0,73,73,128,64,0,0,0,0,136,0,0,64,0,0,73,72,0,346,128,128,64,64,64,0,128,128,64,72,136,128,136,64,64,148,148,148,149,147,157,148,157,156,157,148,156,229,156,229,229,220,221,301,437,293,436,301,438,228,294,294,156,228,367,437,220,156,75,364,74,73,156,147,74,220,219,74,220,229,157,83,147,293,157,220,229,229,228,219,293,439,366,291,445,373,301,365,219,292,292,365,365,228,292,228,229,219,0,0,0,64,137,137,137,136,128,128,72,0,0,0,0,0,0,0,0,0,0,64,64,64,64,64,64,0,145,64,0,0,0,0,0,64,0,64,64,64,128,128,128,128,209,64,64,64,64,72,8,8,219,148,2,148,148,157,75,221,147,147,229,157,74,229,229,229,302,221,436,365,220,438,302,293,229,148,229,293,294,291,219,147,155,211,293,75,302,229,83,147,229,9,73,155,156,9,83,219,165,229,293,157,228,229,220,156,437,292,446,291,364,438,437,502,292,365,220,356,220,292,300,218,128,137,301,147,292,284,147,210,64,64,64,192,200,136,136,64,64,145,200,128,64,64,64,137,72,8,0,64,64,64,64,64,64,64,0,0,0,0,0,0,0,0,64,209,128,64,0,73,136,8,0,72,282,148,157,221,147,148,157,149,293,147,164,229,221,228,302,229,366,302,292,437,301,437,301,365,302,302,294,147,229,291,283,437,437,373,292,75,229,229,74,147,157,229,219,0,229,83,83,73,147,156,229,157,220,293,366,439,446,365,501,438,510,502,511,502,493,429,438,437,365,511,511,292,437,293,228,147,148,220,283,220,284,291,291,200,64,72,0,72,128,200,136,201,72,64,128,128,64,72,137,64,64,0,72,64,64,0,64,64,64,0,0,0,64,137,209,72,0,0,0,64,136,0,72,8,81,73,157,156,157,220,149,157,149,284,156,156,375,229,375,221,367,303,228,365,365,436,373,437,293,366,294,220,365,292,292,301,301,82,364,373,301,229,155,147,157,220,156,220,229,156,74,0,147,84,229,157,220,156,301,364,372,220,429,365,501,365,366,438,510,509,502,374,511,502,300,510,511,429,438,439,293,148,356,365,147,292,292,228,428,355,200,136,0,8,0,64,273,200,0,0,64,73,0,64,209,73,8,0,0,64,64,64,64,64,64,64,64,64,64,0,0,72,64,64,64,0,0,8,8,0,0,221,84,156,220,149,156,149,157,156,366,156,229,156,293,302,228,366,437,364,365,365,229,293,221,294,437,429,436,428,301,436,373,437,365,372,293,301,229,229,148,220,156,229,147,73,146,83,156,229,229,221,229,293,445,292,511,429,501,446,502,437,501,510,511,511,510,509,501,510,437,511,210,437,365,437,365,301,293,147,228,365,364,429,301,283,136,128,136,64,0,0,64,64,0,0,0,0,0,0,128,64,64,0,8,8,0,64,64,64,64,64,64,64,64,64,64,0,0,0,73,136,0,0,72,0,157,84,220,221,157,147,156,156,221,220,229,156,365,302,221,219,365,292,293,439,365,293,229,294,228,365,364,437,371,436,300,427,364,373,300,301,373,228,228,147,147,74,156,221,292,148,74,229,220,157,229,229,228,438,437,501,510,510,510,445,437,501,511,511,510,511,500,509,511,511,365,438,437,437,292,446,365,293,147,292,218,292,429,292,356,208,64,64,128,136,145,72,0,0,72,0,0,0,0,0,0,64,64,64,64,64,0,0,72,72,136,209,136,0,0,0,0,0,0,0,0,0,0,0,64,157,148,83,220,148,83,156,148,284,229,156,293,228,228,228,365,365,293,366,366,228,302,220,220,293,365,301,226,509,510,500,510,435,438,292,436,294,302,83,147,1,148,219,221,221,156,229,157,229,229,157,301,164,365,511,501,429,500,445,509,437,509,501,501,501,501,502,510,437,502,510,502,373,510,429,437,439,293,229,292,283,301,429,292,293,501,346,0,0,128,136,72,8,0,0,0,0,8,0,0,72,73,8,64,128,128,64,64,64,64,64,72,137,0,64,73,0,0,0,0,137,0,0,64,64,157,157,148,221,83,220,219,148,293,156,293,220,229,220,292,437,293,301,439,293,302,366,294,229,292,301,437,500,510,499,417,499,371,437,419,364,366,357,157,73,146,156,148,229,148,156,221,156,156,157,293,511,429,511,438,437,501,509,501,437,503,437,445,436,436,502,446,437,502,437,502,501,510,437,374,292,365,220,147,291,365,293,365,293,292,292,427,281,64,0,136,136,136,72,0,72,0,0,200,136,72,8,0,8,72,0,0,0,136,64,64,64,64,64,64,64,136,0,128,72,64,0,64,64,0,148,221,156,157,148,283,84,292,157,229,292,301,293,437,437,228,301,366,364,302,294,375,229,293,366,437,154,436,510,510,499,511,435,436,373,365,429,148,229,156,157,148,229,157,229,156,156,83,221,156,365,511,366,511,438,510,437,510,445,509,510,509,509,510,510,501,511,446,510,437,510,438,511,511,438,366,292,364,74,429,365,293,510,366,301,292,364,283,145,0,0,136,136,128,9,0,0,0,0,0,0,64,64,0,0,0,0,64,64,64,0,0,0,64,145,273,64,128,64,72,0,64,64,0,0,157,220,220,84,211,149,148,221,229,292,293,293,293,228,437,302,293,293,293,302,366,293,229,366,366,364,292,373,373,364,510,508,354,437,292,309,229,148,156,228,74,157,157,157,156,157,84,157,156,157,511,228,429,301,502,438,510,510,510,501,511,501,509,445,437,511,510,436,437,510,511,437,438,502,365,438,301,356,147,365,364,292,291,293,365,292,292,429,291,218,72,0,136,136,72,0,136,72,72,64,0,73,0,0,0,0,0,0,0,0,0,0,0,64,64,64,64,64,72,73,64,64,64,0,72,156,156,157,148,219,84,293,157,293,156,294,293,220,292,293,302,292,301,294,228,293,229,366,366,438,229,292,436,363,363,373,373,365,509,500,301,148,229,91,292,229,156,221,156,157,157,157,157,156,229,511,365,374,365,510,502,511,509,437,510,510,510,509,509,508,501,437,510,445,511,511,511,374,439,447,374,293,292,294,437,437,366,300,301,365,365,301,501,291,156,219,64,72,136,136,64,64,0,64,64,64,64,64,64,64,136,128,128,64,136,136,136,128,64,64,0,0,0,64,64,64,72,209,128,128,148,220,148,282,156,292,221,221,293,294,294,228,301,293,301,293,301,293,229,293,301,293,367,438,292,156,156,301,436,301,437,436,373,219,364,229,229,83,156,83,293,157,157,148,156,156,157,156,221,301,437,229,438,365,510,501,511,511,373,501,509,509,499,510,499,507,511,438,510,511,445,510,373,511,365,364,365,292,219,364,437,301,365,373,365,292,365,365,292,147,138,147,355,64,128,136,64,72,145,0,0,0,0,0,0,0,64,64,64,64,64,0,0,0,0,64,64,209,0,64,200,128,128,128,128,156,147,282,219,221,293,157,293,220,294,294,292,292,301,293,292,292,301,365,437,301,293,439,229,165,147,229,301,301,501,364,437,156,229,294,229,84,229,91,155,229,148,148,229,229,229,229,228,229,302,502,293,438,437,429,510,501,510,446,510,509,499,498,499,425,499,509,511,510,510,510,510,438,511,438,437,438,293,292,437,365,365,365,365,365,301,365,292,228,83,73,220,210,137,64,64,136,8,0,72,72,0,0,0,0,72,64,64,64,0,72,0,8,64,64,0,64,64,64,128,64,0,0,0,201,148,220,219,220,292,221,221,220,229,302,292,301,365,302,228,420,365,300,293,365,365,366,365,229,148,156,229,147,220,293,156,301,302,229,229,148,164,156,229,301,229,156,157,301,157,229,237,293,229,229,438,438,511,511,375,510,445,510,446,509,511,509,490,490,416,508,508,365,511,510,447,511,438,511,439,502,365,292,293,437,429,437,373,365,437,365,365,292,147,156,73,146,147,201,136,64,64,136,64,218,72,8,73,72,72,72,0,64,0,0,64,128,64,0,0,64,64,128,64,0,0,0,0,0,201,147,219,220,293,293,221,220,229,293,229,292,365,292,302,283,282,364,437,364,293,366,439,292,221,75,74,147,291,75,147,74,148,156,229,148,229,229,156,229,220,220,221,229,157,230,364,365,301,229,293,229,438,439,510,438,510,511,510,502,500,511,510,509,499,426,498,509,511,438,437,437,511,429,511,292,366,374,301,300,508,428,438,365,373,292,365,365,365,83,156,83,155,155,156,219,136,136,136,72,8,209,73,0,0,0,72,8,72,72,72,0,0,0,0,64,128,128,0,0,0,0,0,0,0,0,220,220,283,220,220,221,

293,229,294,228,293,219,228,230,355,293,364,437,300,366,439,365,229,147,74,74,229,65,148,74,155,228,156,148,165,229,365,220,221,356,429,229,230,221,230,230,230,229,229,229,229,438,511,437,510,439,510,511,511,501,437,510,508,510,509,499,510,365,437,510,429,511,429,447,301,374,366,228,354,436,501,228,365,365,292,373,364,365,220,82,228,356,156,83,156,65,136,64,64,72,8,8,64,145,72,72,72,8,8,8,0,64,72,137,136,136,73,64,64,72,145,72,0,0,0,220,147,292,228,221,293,229,228,293,293,292,220,292,303,356,366,437,437,366,374,301,165,147,73,74,156,73,74,74,147,9,221,220,229,229,229,229,293,430,366,366,366,293,221,229,229,230,230,230,230,301,301,446,438,510,510,438,511,510,502,501,445,510,509,509,510,509,502,511,510,501,510,439,301,511,429,229,292,508,437,510,228,365,365,365,365,292,293,293,156,228,301,148,156,219,1,84,137,136,64,64,64,72,0,0,8,8,0,128,128,64,64,136,136,128,128,128,136,64,0,0,64,72,145,73,229,156,293,229,293,293,220,228,228,293,301,293,365,146,365,284,282,366,366,438,292,147,74,147,83,74,64,156,156,156,229,292,302,220,229,221,438,438,430,366,365,293,294,366,301,229,229,229,220,293,293,302,438,438,366,301,439,511,436,511,510,509,501,509,509,509,509,501,511,502,510,510,374,439,374,364,293,428,508,510,364,227,365,365,301,364,301,221,293,156,228,147,156,220,146,75,84,148,216,64,136,136,128,128,64,128,128,128,128,128,136,136,136,128,64,8,0,0,72,0,0,73,73,8,17,293,283,221,229,302,229,219,228,155,302,437,301,293,356,229,292,437,366,366,292,156,75,229,82,156,64,155,220,293,293,293,302,302,293,230,293,365,229,229,156,156,365,439,439,366,293,365,293,230,293,429,374,229,438,511,365,374,511,510,508,510,509,510,510,510,509,509,510,510,438,511,511,438,373,439,229,220,435,363,428,437,501,365,301,301,301,301,228,292,293,229,220,83,228,74,148,83,83,146,65,2,73,75,145,81,145,136,72,73,72,282,136,128,64,64,64,0,0,8,9,9,9,9,9,8,219,292,157,229,294,229,228,220,294,366,437,292,356,428,364,438,437,438,438,301,146,229,73,74,73,219,229,365,294,230,220,156,149,221,293,292,366,366,438,438,375,374,438,366,375,367,367,439,366,294,366,366,301,293,439,511,438,438,510,501,511,501,510,509,509,501,501,510,510,511,502,437,438,438,366,229,293,435,372,510,437,437,364,301,301,300,156,228,292,293,228,292,156,219,147,149,148,138,145,73,74,73,75,146,74,81,137,74,138,282,136,128,128,0,64,64,64,64,72,64,0,8,0,0,0,302,292,156,302,230,229,228,293,293,437,437,292,355,437,364,217,438,365,365,220,147,155,146,74,148,293,302,229,229,156,220,438,292,84,84,84,285,219,366,439,366,439,375,366,157,148,293,438,439,438,294,302,302,156,438,511,511,438,511,447,511,510,437,301,510,438,508,510,502,438,510,438,438,365,302,229,429,508,365,428,501,364,364,228,228,365,229,220,293,156,228,220,228,74,84,76,147,138,146,137,146,81,74,219,74,146,211,74,146,128,64,0,0,0,0,0,0,0,0,8,64,64,8,73,64,303,292,220,302,229,229,228,366,366,436,437,365,364,437,355,437,366,365,301,147,292,146,146,157,429,229,302,293,501,437,293,156,220,220,293,365,438,430,366,438,367,293,438,439,375,293,292,293,292,301,367,294,366,301,438,510,511,439,511,511,437,510,510,510,509,511,509,438,511,437,511,356,438,429,221,365,435,435,437,364,501,428,292,302,301,156,156,229,293,229,301,220,219,74,84,147,147,138,138,137,82,82,73,218,147,74,146,82,65,0,0,136,128,64,0,0,0,0,0,0,0,8,0,0,8,303,229,229,294,302,293,365,302,366,437,437,356,291,437,365,437,366,365,229,156,73,72,148,230,365,302,302,365,220,146,219,365,219,228,229,156,156,220,366,366,366,366,439,302,366,439,439,302,293,357,229,301,365,374,366,438,511,511,510,510,511,510,510,365,437,502,438,510,365,438,511,437,511,366,292,436,499,437,436,365,437,510,365,155,228,229,164,228,293,228,228,220,74,84,157,83,66,210,146,138,146,154,139,219,75,73,73,64,0,64,137,136,209,136,136,128,72,0,0,0,0,0,0,0,0,302,229,229,302,293,357,437,294,366,501,437,355,437,437,365,364,365,366,220,229,219,74,221,156,365,302,220,365,437,293,221,221,221,294,294,294,294,294,294,302,366,374,375,375,366,156,293,375,375,366,293,366,229,229,374,366,294,293,366,429,511,366,438,301,366,366,293,510,447,439,365,438,365,221,436,436,508,436,436,365,502,510,365,155,156,292,229,292,155,293,429,147,75,84,83,84,1,210,138,73,73,154,146,72,76,138,82,137,0,357,137,146,137,64,211,74,128,0,9,0,9,0,0,0,0,302,230,230,302,293,357,438,302,429,500,364,356,365,365,155,365,228,301,220,156,82,156,229,229,366,302,364,365,365,229,366,366,365,365,293,366,365,229,230,294,294,302,302,294,375,366,366,367,365,366,229,229,294,294,229,230,366,158,229,302,502,511,502,438,511,438,292,438,439,511,292,438,229,221,500,363,435,509,364,364,501,300,228,155,221,229,229,293,157,229,155,74,84,84,75,147,65,211,74,74,137,146,83,73,83,74,137,0,146,293,72,219,218,64,74,75,210,137,0,8,73,0,0,0,0,302,293,229,294,293,365,502,365,428,437,355,365,437,229,219,439,228,220,156,220,229,156,229,365,230,294,365,229,228,366,294,366,366,366,229,375,302,229,293,430,429,229,294,230,221,220,302,439,366,430,301,229,293,294,229,293,230,156,293,229,439,219,438,365,237,365,375,447,301,374,374,365,229,228,435,355,501,508,364,364,501,301,228,229,228,229,292,229,165,429,146,75,85,156,84,147,146,220,73,219,146,73,75,73,146,219,73,64,75,220,72,219,282,64,146,74,218,0,64,0,1,0,8,0,0,293,292,229,229,293,293,429,363,290,501,356,365,438,302,294,366,229,147,229,229,83,229,364,220,230,375,302,221,365,501,302,229,148,156,293,292,293,293,229,293,365,438,365,293,294,221,148,228,374,374,439,439,293,294,230,229,302,229,157,230,366,228,301,511,511,293,155,438,375,438,301,365,229,301,436,436,437,508,364,365,437,301,292,301,229,229,301,157,229,228,65,84,84,221,84,147,74,74,209,202,138,73,219,146,64,136,0,146,66,156,0,210,283,64,211,138,137,138,137,136,73,1,0,72,64,229,292,293,229,293,429,502,501,436,291,356,301,301,293,229,293,147,302,229,229,83,294,365,230,302,365,229,365,293,230,293,429,228,365,220,220,148,147,220,229,293,301,373,437,437,366,229,148,148,438,366,302,366,293,293,230,302,302,221,157,221,156,292,293,229,292,155,438,229,365,293,220,302,364,436,437,437,437,437,436,437,365,437,293,228,301,229,164,229,146,83,74,74,75,148,148,74,74,209,73,74,73,73,146,136,64,282,156,74,0,0,219,209,64,64,0,65,0,65,1,73,72,0,9,0,365,228,293,293,292,501,437,437,429,283,356,437,229,294,229,366,156,367,229,229,229,229,229,221,293,365,301,356,293,293,365,293,284,429,356,357,301,365,366,301,293,366,294,220,437,365,365,292,301,220,365,366,302,147,229,294,229,157,294,229,148,221,220,229,229,301,164,293,229,293,293,156,366,292,438,365,364,437,364,501,365,365,365,293,229,300,293,229,229,73,83,75,220,147,147,83,147,147,210,137,74,73,137,136,64,283,210,156,147,229,0,209,73,64,128,64,138,66,82,145,137,136,64,0,8,284,293,294,294,220,429,437,501,438,356,356,365,229,301,229,365,229,230,229,292,229,148,220,438,502,301,220,293,365,155,374,156,229,229,220,156,156,293,292,220,292,293,366,366,229,365,365,293,220,301,365,292,366,302,228,156,294,147,229,294,221,74,221,229,293,156,164,366,301,155,293,229,366,365,437,372,300,438,501,436,365,365,292,229,229,301,156,229,300,146,74,147,147,210,220,147,75,147,74,145,74,74,137,209,155,229,148,155,147,155,1,64,192,328,264,64,65,82,73,18,18,346,136,65,0,284,228,293,292,293,364,365,509,438,355,293,437,229,229,229,293,220,367,229,229,156,221,292,437,365,293,301,301,156,366,229,429,429,439,439,302,157,229,229,293,293,357,292,293,293,156,148,365,365,221,365,301,365,302,294,148,83,293,156,157,302,147,229,302,157,221,229,438,228,221,82,293,229,365,365,436,437,365,436,372,365,292,228,229,229,301,228,228,300,73,147,147,74,211,10,147,147,76,66,138,218,74,210,146,156,220,148,155,212,147,146,201,218,273,328,65,0,73,9,9,73,73,137,128,0,209,219,292,229,365,428,511,373,301,437,156,437,229,220,220,366,293,375,221,293,221,157,291,437,501,437,365,284,365,294,366,301,229,157,157,221,292,293,156,156,156,293,366,365,219,365,293,365,365,366,292,301,365,229,303,294,75,293,147,156,366,229,220,221,157,220,302,294,228,229,74,294,229,300,365,437,364,365,436,365,429,292,302,229,229,365,229,228,292,146,75,74,75,219,147,147,147,75,147,74,217,138,355,210,91,164,219,156,292,220,147,200,328,209,210,65,65,73,73,65,18,9,73,128,128,209,283,228,293,366,501,439,438,365,437,156,437,156,365,220,365,221,294,221,293,221,156,292,221,429,293,364,502,501,429,302,229,221,221,221,221,229,220,366,229,220,293,366,302,365,430,365,366,365,366,366,219,375,293,293,229,293,75,229,147,366,221,147,294,157,156,447,230,294,294,220,365,229,428,437,365,292,365,228,365,365,356,293,293,293,292,293,229,229,138,74,147,74,74,155,75,155,147,74,73,66,217,74,218,155,92,283,220,366,65,65,201,201,265,264,73,0,355,1,10,9,1,73,136,64,137,146,220,293,439,501

,439,366,365,429,156,429,301,229,365,301,220,293,229,229,293,220,156,157,501,293,229,230,365,366,366,365,429,430,229,156,229,229,229,229,375,293,293,365,292,365,429,365,366,365,294,221,365,375,294,375,229,74,157,148,293,219,293,365,229,229,511,229,429,302,365,293,293,364,502,364,437,365,438,437,292,220,229,229,147,292,301,292,229,74,74,147,75,74,147,147,148,283,147,146,74,74,146,291,155,155,283,219,283,83,137,264,274,210,264,138,74,138,64,73,9,146,145,72,210,74,156,292,293,439,284,366,365,438,429,292,365,437,301,292,302,293,292,229,230,229,292,147,294,148,501,229,228,365,510,511,511,439,365,365,292,293,83,83,156,221,230,229,229,365,364,292,365,365,375,365,294,365,366,302,293,367,293,221,83,366,147,9,220,229,365,438,367,429,511,365,294,374,510,437,365,437,227,510,437,365,229,293,229,155,365,429,229,228,138,146,74,83,74,147,219,76,148,155,82,147,218,218,210,82,164,282,219,356,221,138,264,137,65,74,73,1,209,74,9,0,0,73,64,137,147,220,292,293,374,293,439,366,439,220,355,365,501,365,221,301,292,284,229,294,147,357,139,148,366,366,438,229,229,301,365,500,438,366,365,365,156,157,148,83,83,147,148,229,365,293,365,292,365,429,366,437,229,301,365,365,366,302,229,220,366,147,219,156,220,430,302,294,439,374,293,221,292,510,373,437,364,364,365,429,301,301,229,429,148,501,357,301,220,220,73,2,74,147,147,147,76,83,219,221,74,74,217,146,73,156,282,147,356,148,1,1,65,65,0,73,1,146,0,73,72,81,64,1,8,156,138,292,220,439,230,439,302,447,429,209,356,500,293,365,437,365,211,229,367,302,301,294,284,229,293,302,366,229,229,293,438,366,293,301,373,366,437,365,156,156,74,75,75,293,365,303,293,365,365,429,365,302,301,366,366,293,294,366,220,439,293,139,302,221,220,293,221,302,156,229,157,501,429,301,429,438,437,502,364,229,302,292,364,292,356,157,301,229,293,73,73,2,138,147,75,220,229,219,438,82,157,146,145,145,76,217,211,283,147,137,146,65,73,282,65,1,65,65,65,0,154,1,81,145,229,346,429,156,438,366,438,294,439,437,502,356,501,229,219,293,293,147,221,293,294,228,294,221,375,375,157,293,438,438,293,365,439,439,366,229,301,156,366,365,229,293,292,75,83,147,229,366,365,301,301,293,229,302,366,374,365,438,302,301,366,447,148,229,156,227,229,220,302,228,229,229,436,365,301,501,364,501,502,292,229,229,229,292,365,366,84,374,301,293,156,73,73,74,74,147,146,145,155,155,365,301,82,74,138,148,218,74,155,146,137,292,137,64,73,73,138,137,0,0,0,154,137,81,64,156,355,292,293,439,439,502,365,439,292,429,364,428,229,293,293,294,220,220,157,229,366,293,294,148,301,375,84,293,366,374,229,219,438,374,302,302,229,84,366,374,302,230,293,83,83,147,293,366,365,156,229,301,302,302,366,366,438,302,301,366,302,157,293,220,365,229,229,302,229,230,302,436,365,302,364,429,510,438,156,301,302,301,365,292,293,83,438,293,293,220,155,74,75,138,147,219,157,82,82,365,148,74,146,145,148,356,74,155,0,128,220,138,72,209,289,281,280,64,64,0,0,81,73,137,74,356,284,365,356,366,284,430,503,220,365,282,364,293,294,302,147,230,293,157,157,294,302,293,302,148,149,374,366,229,229,229,229,220,366,429,430,366,229,156,301,228,294,230,229,156,148,220,367,229,229,156,301,301,157,439,366,438,375,220,439,156,439,365,147,294,230,428,229,228,293,228,510,374,301,364,365,510,365,228,365,293,300,373,293,156,83,366,438,292,502,229,147,148,74,293,220,91,146,373,91,373,155,83,146,220,219,147,155,217,64,220,137,64,64,288,426,425,128,0,74,9,154,73,72,292,292,356,212,430,430,439,430,447,229,429,364,356,356,365,228,229,75,230,357,157,294,293,367,230,230,293,85,221,157,157,293,302,229,156,84,293,228,365,302,229,221,220,293,229,293,147,220,229,293,302,301,367,365,156,302,302,229,375,221,438,302,511,366,229,147,230,365,221,292,302,219,510,438,364,372,301,365,292,293,364,364,365,437,293,156,83,301,292,301,365,220,293,75,138,365,293,220,91,154,292,227,374,82,145,147,218,147,219,281,136,137,64,64,0,209,272,344,136,73,73,74,73,73,64,221,293,356,219,365,229,439,447,439,437,365,365,293,356,293,229,302,147,229,292,220,229,229,229,294,230,229,293,230,294,365,430,365,438,365,365,228,147,221,366,302,148,230,220,229,229,293,228,439,293,293,292,303,373,301,230,220,155,148,148,220,439,374,375,157,147,230,229,229,301,229,292,501,510,509,373,365,435,301,365,364,300,364,437,302,220,156,220,228,301,365,292,228,147,74,292,147,156,83,155,292,228,90,82,73,218,281,65,147,138,73,73,73,210,64,146,138,138,73,73,81,82,74,73,10,285,293,356,74,429,439,438,439,438,438,293,292,438,438,220,365,294,366,284,294,365,229,222,230,229,366,229,230,229,302,229,229,148,75,75,139,220,301,365,156,229,302,156,229,147,156,148,293,229,293,365,229,229,302,301,157,229,365,220,156,293,301,221,302,366,229,230,229,229,229,230,302,364,510,435,365,437,363,301,429,292,365,437,364,293,228,220,229,228,229,365,301,147,74,75,220,148,147,157,145,227,82,365,155,146,219,292,65,146,202,364,292,291,219,356,356,356,291,291,0,145,145,82,73,73,148,293,291,73,430,365,365,284,438,439,293,357,365,366,229,365,365,366,292,229,293,357,229,230,229,293,366,366,294,229,366,156,156,293,220,366,293,148,156,301,220,229,302,147,156,148,156,230,357,221,302,229,301,367,301,302,293,366,147,221,229,294,221,294,302,221,230,230,229,229,230,220,365,501,435,301,435,364,365,301,292,437,510,293,229,228,293,228,365,292,156,301,139,74,219,147,220,148,145,145,291,301,155,82,146,219,219,74,147,283,365,292,282,283,64,210,218,210,145,65,218,73,82,281,137,148,292,292,146,292,429,293,365,293,365,293,293,293,438,365,501,301,292,438,221,83,220,220,439,156,367,230,230,229,293,366,294,294,302,365,157,294,229,156,156,301,302,365,294,148,157,147,156,301,221,302,293,301,292,302,374,302,294,229,220,221,221,439,293,293,230,230,230,230,230,293,364,373,502,435,301,362,365,428,292,437,437,364,229,366,220,228,301,365,293,83,228,75,75,292,76,147,148,145,146,292,301,82,73,74,283,146,73,147,218,364,356,283,64,128,128,72,65,74,65,73,74,73,208,137,220,364,284,220,229,220,293,429,229,302,366,229,292,503,366,219,365,220,365,430,293,75,229,293,157,294,229,302,230,293,301,157,157,293,229,294,294,230,229,157,221,366,365,366,293,148,156,74,293,293,229,302,447,366,302,374,301,293,220,73,220,221,374,302,221,231,293,230,301,229,293,437,373,437,436,365,500,364,501,365,437,437,221,229,293,156,301,237,365,148,156,220,75,75,147,220,147,148,145,145,293,227,83,155,146,228,74,73,219,283,364,292,136,137,283,283,355,146,73,65,145,9,1,1,219,147,221,220,140,437,293,228,293,293,229,429,229,365,365,430,156,156,302,84,292,365,293,76,156,365,293,221,230,367,302,375,303,294,229,230,148,230,293,430,157,148,156,293,229,292,220,148,219,220,293,229,302,438,293,229,438,301,292,228,293,156,294,366,221,365,439,365,228,366,229,302,438,502,510,364,510,500,356,364,365,437,292,229,228,229,229,365,374,147,229,156,147,74,219,76,357,147,146,145,145,300,91,292,146,90,356,147,282,283,138,136,136,283,218,283,291,218,210,1,81,73,154,282,209,364,212,148,356,148,292,293,438,221,220,502,365,365,229,438,511,366,156,366,229,84,219,366,230,157,148,285,228,429,366,366,438,366,367,230,157,230,294,375,364,366,84,229,366,293,221,438,147,147,211,229,229,302,437,302,157,364,301,438,293,228,221,230,367,148,221,229,302,294,302,229,229,438,219,429,301,511,436,365,364,510,501,220,228,373,220,293,301,365,83,301,293,74,75,219,148,228,147,145,145,211,146,73,147,147,229,293,292,74,138,128,346,283,219,73,73,65,64,0,64,72,9,209,73,209,282,221,221,212,156,75,293,365,292,229,293,220,502,156,83,511,438,293,439,366,229,84,147,301,302,230,230,221,148,156,148,367,375,230,158,157,230,293,375,293,439,285,220,366,293,366,374,365,74,147,229,437,438,437,366,293,227,301,438,293,156,149,293,148,221,229,156,365,366,374,302,293,293,220,438,365,428,364,501,438,437,292,220,229,293,228,228,438,366,147,365,220,74,148,156,149,156,147,146,219,148,146,292,219,229,146,146,354,219,146,65,137,283,210,137,128,64,0,0,64,73,8,146,146,209,291,221,229,149,355,220,357,293,365,229,293,365,293,230,220,438,502,502,366,439,366,294,221,220,365,293,375,294,229,221,230,229,156,220,293,375,439,438,293,220,439,365,221,375,357,367,228,293,147,147,148,365,365,301,374,301,365,301,365,229,156,149,302,148,375,229,229,293,302,165,229,301,229,229,228,293,429,292,428,292,365,437,237,301,221,293,229,365,156,220,228,75,74,220,156,148,157,84,146,149,146,145,82,146,84,156,82,219,146,293,292,138,64,218,282,355,209,137,137,64,137,82,138,146,210,356,293,221,293,292,355,364,302,439,430,220,302,365,438,156,148,429,501,366,367,366,365,366,294,74,155,292,366,302,301,366,366,438,366,366,365,293,156,157,229,365,429,221,302,502,294,221,293,220,147,220,365,438,438,366,437,365,366,365,220,156,157,293,294,230,221,302,302,294,165,229,229,229,229,229,365,437,373,501,429,365,438,229,301,229,365,156,301,365,228,147,74,148,219,148,156,284,148,147,158,145,220,147,146,293,83,138,73,210,73,220,293,292,73,64,137,292,291,292,65,73,137,137,146,209,291,220,220,220,219,364

,364,219,375,294,220,293,365,229,302,156,229,357,374,302,294,437,438,438,293,156,83,156,156,220,155,302,293,221,148,220,366,439,229,293,293,366,293,294,439,229,294,293,221,284,220,365,365,364,439,438,365,293,221,156,156,221,221,229,302,230,220,229,302,221,301,301,229,229,293,364,301,365,436,300,437,365,292,156,301,228,156,156,374,365,66,74,292,211,221,220,292,156,219,147,155,148,292,155,220,73,147,73,293,146,73,219,293,292,146,0,64,136,136,273,209,0,74,137,283,291,221,221,220,293,292,356,293,293,439,365,229,149,438,302,229,157,157,293,439,367,229,438,375,221,365,438,365,229,301,157,157,366,229,365,366,375,366,294,156,366,375,293,293,367,220,293,156,229,221,229,365,229,218,365,437,366,229,221,221,157,302,157,230,157,365,157,229,155,229,228,229,156,301,365,438,374,437,436,365,510,438,75,220,437,156,301,156,293,146,75,148,147,148,293,147,147,219,219,147,156,219,219,156,156,228,82,74,147,83,146,136,211,219,146,137,64,75,75,75,1,73,73,65,291,291,148,157,156,220,293,365,439,293,439,438,293,156,293,302,366,293,157,221,293,374,439,301,293,430,302,230,229,220,365,293,229,366,302,221,229,439,438,366,229,302,438,293,229,366,365,229,220,229,220,293,365,229,293,366,302,302,294,221,229,221,357,294,294,302,156,155,293,157,228,219,156,228,365,437,365,510,300,437,437,438,292,75,365,292,229,365,156,364,74,75,293,148,220,149,220,149,292,148,147,156,219,221,83,83,229,9,145,137,155,147,73,146,146,220,291,146,219,292,292,292,147,137,146,291,283,220,148,220,212,293,503,366,229,302,439,293,220,157,294,302,293,366,221,293,229,293,438,365,221,148,156,293,366,301,375,367,375,439,439,438,438,302,302,365,302,301,301,293,366,438,221,228,293,293,293,229,293,356,365,365,156,157,284,221,229,293,229,437,302,156,228,220,157,228,228,156,301,365,438,437,510,365,437,428,437,365,438,437,147,373,147,293,146,75,147,220,292,157,156,148,156,220,148,219,155,292,83,146,74,73,73,73,137,145,145,137,219,293,293,292,283,219,292,293,301,74,137,65,283,281,221,148,75,221,147,293,438,294,302,439,294,301,156,229,302,302,229,156,293,375,303,220,438,438,502,301,301,302,229,438,366,365,229,156,157,375,375,375,366,293,365,293,294,293,438,221,221,229,365,293,293,229,365,293,429,155,221,221,220,221,148,230,437,229,229,228,165,229,155,228,301,373,502,437,501,438,437,364,437,364,365,292,291,292,365,220,284,74,147,219,147,220,147,84,148,220,147,146,146,147,146,73,219,220,293,292,138,218,154,81,292,292,292,293,292,210,73,145,146,146,73,65,138,144,64,220,157,148,157,148,294,365,439,229,366,439,221,293,229,293,229,229,220,156,157,229,366,365,301,365,366,375,302,367,375,375,366,437,437,373,366,367,375,430,437,302,430,302,364,365,221,221,229,293,156,229,365,365,301,301,155,229,302,84,429,157,365,229,301,292,156,229,237,229,293,301,300,438,436,501,373,437,364,437,364,365,220,292,364,147,74,73,283,146,292,292,292,292,292,292,293,293,356,293,365,293,365,365,293,301,218,74,136,136,146,356,365,364,137,65,147,74,147,147,138,64,64,137,64,201,220,148,220,157,147,365,293,366,439,284,366,229,293,229,366,229,229,157,83,292,293,157,156,156,229,229,220,438,438,374,366,229,229,293,293,366,365,293,365,375,366,375,365,366,229,221,229,429,293,229,293,438,229,293,438,148,221,431,158,365,294,155,156,229,156,229,229,228,229,430,301,437,437,427,502,373,438,365,292,220,292,147,438,438,221,146,147,148,219,146,148,146,210,74,147,147,74,138,146,146,219,219,219,292,292,137,74,136,136,137,64,64,64,73,64,0,0,0,283,283,65,64,64,283,274,147,148,148,221,147,221,293,293,439,293,365,229,230,365,293,302,229,156,157,221,147,429,438,293,148,156,229,228,293,367,375,375,366,365,365,439,367,366,375,367,301,293,374,293,147,221,293,293,293,293,293,301,157,365,293,229,221,228,366,156,220,83,156,83,83,156,228,429,221,302,373,436,437,435,373,437,437,438,75,229,301,292,437,147,293,74,147,148,147,148,147,292,149,155,149,220,148,146,146,147,146,211,146,146,219,146,65,137,64,0,73,146,64,73,0,0,64,0,146,283,64,273,283,274,274,148,293,157,149,156,212,293,156,293,366,365,293,230,366,365,221,301,293,156,156,294,375,293,293,501,429,156,220,366,437,438,438,365,365,365,365,366,375,366,366,156,366,438,302,147,221,429,293,293,229,429,301,229,374,293,294,221,302,365,229,220,147,156,156,156,83,155,221,302,293,437,437,373,436,436,437,445,83,220,219,292,510,365,156,138,139,84,84,220,74,220,149,148,148,220,148,219,146,73,147,74,293,82,155,300,228,73,209,73,73,65,65,210,211,147,211,146,74,74,74,137,145,283,282,209,220,221,148,221,147,212,293,366,148,439,438,511,301,373,438,229,156,228,229,229,220,293,229,294,302,293,228,501,501,501,430,365,438,438,366,366,438,293,367,156,301,365,229,429,147,229,229,301,293,437,293,229,374,292,229,157,155,374,220,229,82,156,157,156,220,148,293,229,429,373,437,438,502,437,510,293,373,156,220,74,147,365,220,156,66,2,147,229,147,147,284,148,219,149,220,156,146,146,73,75,439,146,146,365,292,154,365,147,209,210,218,218,65,1,73,211,219,147,146,137,65,145,210,347,209,221,229,294,156,212,148,221,293,438,365,439,439,366,220,439,366,229,293,156,229,229,220,365,293,366,438,438,438,366,302,230,302,302,375,438,229,302,375,156,229,438,366,438,293,148,157,293,301,429,293,293,157,365,229,293,293,366,220,229,293,229,229,82,229,156,292,147,219,365,437,373,373,437,436,438,437,220,229,148,292,156,220,301,75,147,84,148,156,148,219,148,220,148,156,149,147,148,211,73,76,365,365,155,229,155,365,219,74,147,74,74,65,73,64,65,137,219,210,283,209,137,145,209,145,209,293,292,229,302,220,83,220,221,292,439,375,439,439,366,221,293,439,438,293,74,83,156,229,293,430,439,302,293,293,438,439,439,439,366,229,438,374,301,365,220,293,302,366,293,229,221,301,300,429,366,229,228,301,229,221,292,294,374,301,229,237,82,156,365,220,228,156,365,429,438,301,373,437,437,502,437,229,156,301,292,156,365,293,74,212,147,148,220,219,155,211,220,219,156,148,221,147,138,74,76,366,228,219,301,74,155,155,83,139,83,82,64,210,72,0,65,65,1,1,0,64,81,137,145,210,366,356,148,148,284,293,83,229,229,293,439,293,229,366,366,220,365,439,439,302,148,220,147,157,156,156,220,229,293,429,438,366,439,439,439,364,301,365,148,156,293,156,367,221,221,293,301,355,292,228,301,301,229,157,221,366,366,302,365,238,301,156,228,293,220,229,228,219,228,301,373,437,438,510,510,446,220,148,437,220,293,302,292,65,293,219,147,211,84,148,219,219,148,148,220,148,220,139,147,148,292,301,83,292,220,229,73,1,138,83,74,65,293,283,147,140,221,66,65,65,137,145,137,137,137,365,228,147,230,356,220,156,148,221,229,157,293,366,221,366,366,365,365,438,365,366,148,157,157,229,365,293,229,294,375,438,293,229,293,301,302,302,229,156,220,148,220,367,429,301,228,300,365,365,366,301,229,229,148,294,294,302,228,229,228,156,165,365,229,302,220,229,82,229,237,364,437,301,502,502,438,292,301,437,229,220,228,138,65,211,148,82,148,76,147,155,156,156,220,220,155,220,139,147,147,293,229,83,217,147,155,9,9,147,147,74,64,220,218,219,76,221,65,64,65,73,146,210,137,209,293,366,147,220,229,156,147,148,147,156,293,221,221,367,158,293,229,293,356,293,429,147,156,148,148,147,220,221,293,438,365,366,366,438,438,439,366,147,148,221,230,366,366,301,301,228,428,365,229,365,301,229,157,148,302,301,157,156,156,365,156,229,293,229,301,221,147,228,229,301,502,437,437,438,502,301,365,365,148,221,229,301,74,140,146,74,148,220,84,292,76,147,147,156,148,219,148,138,147,83,228,219,83,146,147,293,73,138,65,138,73,65,220,219,219,148,220,73,137,138,146,145,210,210,137,292,366,221,147,221,293,229,74,147,292,156,292,157,438,439,439,430,83,158,293,365,293,357,156,83,83,83,147,148,367,439,302,365,366,301,293,147,156,221,156,229,229,302,228,301,292,291,437,365,301,301,157,365,229,229,157,156,220,229,156,156,229,301,302,229,229,220,229,302,229,373,365,502,438,437,373,437,365,293,292,229,219,65,76,147,155,148,76,219,220,83,146,147,75,147,147,146,138,147,156,228,219,155,228,148,155,138,155,83,138,65,65,219,209,283,292,73,0,0,64,292,218,210,64,64,428,293,221,156,148,221,147,147,147,147,220,220,219,229,228,375,367,430,365,221,366,366,293,229,229,221,156,147,74,83,147,156,221,147,220,147,367,367,148,294,293,366,375,300,293,356,438,229,301,301,157,230,293,158,229,230,156,237,157,220,221,220,82,229,229,292,229,301,229,229,436,365,437,291,373,437,365,293,373,228,229,74,74,146,211,146,147,219,220,148,147,75,147,66,147,82,138,146,76,156,229,156,156,156,155,301,228,156,156,1,1,0,138,219,137,291,137,0,0,81,291,210,65,65,65,364,156,230,294,220,75,147,156,148,75,148,219,220,365,219,302,365,302,366,293,365,438,429,229,83,156,221,220,156,156,221,229,220,156,221,366,156,148,148,302,365,367,220,302,292,355,511,302,364,301,221,293,230,229,229,229,302,229,230,156,229,293,220,220,229,228,293,292,302,300,290,301,365,301,437,292,373,220,364,229,301,138,139,74,83,147,148,147,292,283,82,82,76,146,75,147,74,73,148,220,228,164,164,155,293,293,155,147,1,146,82,65,1,0,64,64,73,0,64,64,137,1,0,73,137,220,148,229,230,

156,229,292,219,220,221,84,147,219,75,156,229,83,365,301,228,357,293,292,366,365,157,148,294,302,366,229,156,148,83,147,366,294,157,365,365,366,229,147,374,356,355,229,374,428,293,366,294,301,220,302,229,302,229,374,220,293,156,156,156,293,156,301,365,292,293,373,365,292,365,300,365,437,301,365,229,356,65,147,148,219,148,220,147,147,155,147,146,74,155,146,211,74,75,147,220,147,229,148,155,227,82,147,155,82,146,229,228,156,83,82,64,0,0,0,64,0,73,73,65,65,158,284,147,149,147,82,83,220,220,147,155,75,147,148,149,74,147,229,83,156,157,157,157,157,149,156,74,82,83,82,74,82,82,155,293,220,294,429,302,294,301,302,236,437,356,292,302,366,293,430,221,294,229,301,230,293,366,366,293,156,302,293,364,165,292,365,156,365,437,291,373,438,365,438,510,437,437,292,301,301,146,74,139,147,84,219,212,147,155,147,218,75,219,220,147,147,65,148,148,220,219,283,91,146,147,82,228,83,219,156,219,83,301,1,146,137,65,0,64,0,65,137,138,74,1,229,230,147,229,229,220,155,83,147,147,74,74,83,156,156,84,149,74,229,229,156,156,156,157,157,157,157,148,83,82,74,74,73,74,74,156,229,294,156,365,282,302,220,428,355,293,294,356,221,220,294,293,294,221,156,220,221,157,229,229,365,365,229,292,511,293,292,365,290,437,374,373,373,365,365,437,437,365,229,365,138,212,75,356,75,148,148,146,219,283,155,356,147,146,147,146,74,83,148,219,356,364,83,163,74,74,164,155,293,228,74,219,75,82,74,73,0,64,137,137,146,0,0,65,73,229,221,149,228,220,155,148,228,220,220,147,83,84,84,146,148,156,84,148,148,221,230,229,85,149,149,221,220,220,74,74,74,74,220,229,229,294,302,156,355,293,300,302,355,438,293,366,147,221,293,293,229,366,157,438,438,438,438,438,366,221,229,293,366,302,366,300,374,365,291,438,373,365,373,429,437,301,365,301,364,73,148,147,147,211,147,76,147,211,219,147,146,83,210,211,65,147,76,219,212,364,356,164,73,228,147,147,83,229,82,147,82,83,73,73,146,0,137,65,0,65,1,0,65,1,229,220,158,229,155,147,157,219,155,292,220,146,147,83,75,74,74,148,156,83,221,221,148,229,294,293,229,230,229,230,157,221,293,220,294,229,230,294,156,220,438,366,439,511,438,229,228,156,294,229,301,293,156,501,365,365,293,293,229,293,439,302,302,375,375,365,374,438,438,365,437,437,365,437,365,437,502,293,292,283,138,139,291,75,284,147,73,148,283,147,75,74,148,146,283,74,220,76,219,212,356,220,155,155,74,138,210,146,155,82,146,155,73,65,1,0,65,64,0,65,0,0,65,0,73,221,82,149,220,220,220,157,222,219,138,219,221,75,148,148,156,147,83,148,83,147,83,148,148,148,148,83,148,156,157,221,229,229,230,221,156,230,220,221,302,438,366,439,439,301,294,293,156,302,302,228,229,365,437,293,430,365,438,366,439,157,357,301,302,365,292,364,293,372,437,437,438,373,437,300,301,437,301,365,211,138,292,211,147,220,147,211,147,147,76,75,76,84,138,73,74,148,220,284,76,356,219,91,220,228,74,146,211,83,83,356,220,137,73,73,73,0,0,73,74,1,1,1,65,73,157,73,147,156,219,138,228,149,158,147,74,147,292,148,220,220,230,156,156,147,157,157,157,157,220,156,157,148,157,157,147,229,229,229,220,229,294,355,293,294,437,438,447,511,437,429,365,221,302,293,301,229,438,430,365,365,365,301,220,149,366,357,294,293,292,301,437,301,437,501,510,511,437,365,373,301,365,438,301,146,138,146,147,219,219,66,149,211,74,147,212,75,156,147,73,220,148,292,148,139,291,210,82,74,74,2,146,292,83,83,220,210,73,73,83,73,64,0,138,65,0,73,73,65,137,75,212,74,220,220,147,147,292,157,228,228,301,366,156,221,292,228,220,149,84,156,83,156,157,157,157,156,147,292,157,294,292,157,228,220,229,293,355,220,293,501,438,374,511,365,438,365,221,293,292,428,228,302,428,437,157,149,157,302,430,293,366,439,292,221,229,365,229,437,437,510,437,437,437,373,301,365,437,293,138,219,138,138,283,210,147,146,138,147,75,147,76,147,65,211,220,84,147,148,210,148,218,155,155,74,74,219,292,148,228,74,293,138,138,138,137,73,0,64,137,1,0,1,73,146,147,147,73,147,221,221,156,147,220,221,229,302,356,228,291,363,291,292,229,156,156,157,229,157,157,157,157,156,230,147,157,156,83,228,229,293,157,355,210,301,437,366,366,220,293,293,220,220,229,293,294,365,301,365,294,365,438,292,157,229,429,365,366,293,156,302,229,294,501,510,437,502,437,365,438,301,438,438,365,138,283,73,74,283,138,147,147,147,74,147,75,284,73,65,220,220,221,75,76,145,220,217,156,74,74,138,146,147,74,228,74,155,65,0,0,137,0,146,65,138,0,0,146,73,73,156,294,147,148,148,221,157,220,83,293,301,292,364,371,363,355,219,292,365,220,228,156,165,229,156,220,157,156,157,229,148,230,147,229,221,293,221,291,346,438,365,366,439,365,293,301,220,221,221,220,229,301,365,366,293,229,365,157,302,156,293,365,438,366,356,229,293,229,438,510,509,438,373,373,374,301,501,301,429,138,146,73,147,147,74,146,283,75,74,75,147,147,138,138,220,213,293,147,76,146,148,217,220,228,65,146,147,147,218,146,74,73,73,81,146,65,146,282,137,74,0,0,65,65,73,147,146,229,220,221,221,157,229,365,364,365,364,363,363,364,437,438,426,363,291,301,228,292,229,229,156,156,156,83,156,156,155,292,294,229,229,157,292,355,429,228,439,430,211,156,366,220,147,221,220,294,294,230,229,294,229,293,293,293,229,157,365,366,366,365,157,220,220,501,510,501,510,437,437,301,229,438,293,365,146,210,137,147,138,74,146,210,138,138,74,147,73,74,220,220,148,75,211,75,74,219,292,82,155,65,73,148,148,219,284,147,73,72,65,1,354,280,208,137,2,73,137,137,73,73,83,147,75,148,219,294,221,292,292,292,364,428,437,438,366,355,353,437,291,300,362,292,365,292,294,157,156,230,148,147,229,147,220,229,228,228,221,284,347,364,220,510,366,74,366,366,293,229,221,229,221,366,230,157,230,293,157,230,230,367,156,229,366,366,293,220,148,147,502,501,510,510,373,365,301,301,373,301,373,146,138,73,147,74,210,146,138,146,138,146,74,146,74,148,148,219,147,220,75,74,290,82,156,0,64,137,148,148,210,155,292,1,73,65,0,355,418,344,64,66,74,136,137,137,137,156,148,157,74,221,220,366,220,436,363,438,428,363,427,427,365,438,291,292,364,302,228,301,293,229,294,83,229,221,292,229,148,220,155,229,220,157,365,355,355,156,511,438,292,220,293,292,229,221,355,347,292,229,229,230,156,230,230,294,375,229,229,438,366,366,356,157,228,438,501,437,437,437,293,293,365,366,365,301,292,138,73,147,74,73,147,138,138,74,146,138,138,75,293,221,76,220,147,147,210,146,156,291,155,137,64,220,219,210,156,219,210,81,73,65,73,136,274,65,1,139,137,0,0,65,148,220,221,222,221,220,229,293,445,365,217,364,363,364,437,438,437,437,300,365,362,218,301,229,228,294,156,294,230,228,294,156,228,293,229,293,157,355,282,282,220,365,502,438,156,293,439,147,229,283,229,220,357,229,229,221,293,229,292,229,294,293,437,366,366,356,157,293,293,509,502,437,301,293,301,437,365,365,301,364,74,74,147,74,138,74,138,73,74,138,137,74,85,293,149,140,284,140,210,217,228,155,155,72,0,209,148,147,210,155,228,147,82,146,0,1,73,137,73,0,74,64,64,0,65,147,148,148,156,83,148,221,293,365,364,291,428,437,365,438,436,437,437,292,291,355,438,292,229,302,229,222,294,221,157,367,220,229,365,156,293,220,282,210,282,437,219,366,437,219,220,284,220,147,221,283,220,221,221,355,347,292,293,293,229,294,365,292,357,357,293,147,292,438,437,510,373,374,301,229,365,438,301,293,365,138,74,138,147,65,66,74,64,74,137,74,75,220,221,76,148,220,148,356,218,83,147,82,146,146,0,217,146,146,155,146,73,65,74,1,74,73,137,74,0,0,64,73,64,137,74,220,148,157,229,148,228,293,365,291,429,293,502,429,426,509,500,427,436,292,292,299,300,302,294,366,230,156,221,221,366,221,229,302,230,293,293,282,137,221,364,438,220,365,293,365,220,293,84,148,220,292,220,220,157,221,220,284,230,230,437,365,293,229,439,220,147,147,365,365,509,300,365,365,229,365,437,229,502,365,291,74,74,147,74,210,65,73,73,73,75,85,284,76,76,220,75,82,73,82,147,83,155,82,65,65,145,146,147,83,74,137,73,74,73,146,83,210,74,0,0,64,137,65,83,147,157,156,156,148,220,228,293,438,301,293,301,437,437,509,508,490,426,437,365,364,301,300,301,294,293,229,221,229,156,293,221,229,228,230,229,221,211,201,157,364,438,439,229,366,156,430,147,220,156,148,220,437,364,437,429,293,294,221,293,365,365,365,156,439,211,221,229,365,365,502,437,437,293,293,437,357,301,510,365,438,74,74,74,73,137,65,73,73,75,85,219,148,84,219,76,82,146,73,81,147,220,82,73,64,73,145,210,138,220,219,64,73,74,82,82,82,218,65,0,1,64,137,65,74,147,220,156,148,83,220,229,293,365,292,365,363,428,438,509,498,499,426,437,365,437,301,364,293,229,366,229,221,229,221,229,293,229,220,229,294,221,156,428,220,221,365,502,365,229,365,220,156,83,156,156,148,156,229,157,229,367,366,157,229,293,293,356,366,365,220,293,229,365,509,373,437,292,293,373,365,365,429,364,365,220,147,74,74,74,65,65,65,74,84,293,75,147,293,147,283,74,73,73,73,145,82,292,65,1,64,1,210,74,1,1,64,74,220,82,73,82,210,74,0,0,0,65,1,74,148,221,157,

148,221,148,229,374,301,291,437,364,428,502,502,501,501,501,430,292,374,365,365,293,220,229,149,148,157,221,221,221,221,219,228,221,221,220,156,136,157,430,366,438,365,220,156,148,221,147,147,155,220,428,437,366,357,365,301,365,229,356,283,430,357,284,228,292,429,437,365,437,301,293,438,437,293,437,300,292,148,147,138,74,74,73,65,137,76,220,148,148,220,212,219,146,146,73,73,74,73,82,145,74,82,1,82,73,147,147,73,137,74,82,146,75,220,210,146,0,0,0,74,64,82,75,156,148,221,149,293,292,365,365,292,291,365,429,364,500,501,437,365,301,438,365,510,365,229,220,229,148,221,229,220,157,221,74,294,292,230,147,220,221,355,148,221,439,438,430,293,220,156,148,302,293,229,229,293,294,438,429,301,301,156,229,283,292,429,430,228,293,229,365,373,373,437,293,365,292,301,365,365,292,365,76,220,147,73,73,137,137,75,76,76,148,219,148,147,292,219,82,82,74,81,74,220,74,155,73,0,0,64,146,146,1,1,64,0,0,0,0,0,1,0,0,0,82,64,146,148,83,147,285,148,229,220,229,365,292,365,363,292,364,438,437,365,437,438,301,437,438,293,301,156,229,356,220,302,221,220,229,146,229,220,230,147,156,293,229,282,157,219,429,366,293,293,430,292,148,293,293,365,366,366,501,365,229,156,363,355,220,357,293,219,220,228,220,365,437,437,437,219,437,301,228,365,220,292,219,148,292,211,147,73,64,65,76,212,148,83,76,147,292,438,73,219,74,81,81,145,211,83,218,155,73,73,73,147,74,146,361,280,137,65,0,0,0,1,0,0,0,0,73,146,156,83,221,148,148,157,156,228,228,293,438,219,364,363,363,356,364,428,364,293,292,366,293,229,301,221,221,367,302,293,221,157,146,221,228,229,148,292,155,301,219,147,148,365,438,219,366,229,430,302,292,283,355,355,283,292,283,283,347,283,220,292,356,220,292,292,292,220,365,365,437,437,437,300,292,292,365,229,300,211,148,219,220,210,147,73,74,148,148,76,148,148,147,75,364,76,219,82,81,81,82,147,155,219,82,65,64,73,64,74,138,427,200,284,65,292,73,73,282,137,74,64,273,146,73,83,147,84,84,148,148,228,148,292,301,301,229,292,429,365,366,365,437,365,364,365,293,292,157,293,221,294,229,294,84,294,221,74,228,147,229,220,147,156,220,229,365,75,157,293,366,430,365,293,293,366,301,220,156,220,219,283,347,283,284,292,356,284,356,229,292,293,229,365,228,364,292,437,293,292,437,301,292,428,220,147,220,220,211,219,73,76,147,76,147,219,147,84,155,218,364,147,82,81,81,81,145,228,82,73,9,73,0,0,73,146,281,289,210,74,292,137,0,64,0,0,0,9,146,73,74,75,74,83,84,157,157,157,220,220,293,365,229,148,229,301,365,364,301,301,294,229,293,156,294,294,294,222,302,74,302,366,220,292,229,229,219,148,294,220,220,228,227,219,293,357,229,366,293,366,302,292,293,229,229,220,156,220,292,429,283,219,284,430,156,220,357,301,437,365,437,502,437,301,292,356,292,300,292,156,147,220,220,147,147,74,138,76,147,155,156,148,155,219,292,438,147,82,146,136,145,145,300,146,227,82,0,0,74,138,146,137,1,138,138,292,146,64,210,283,283,138,65,82,82,83,148,148,221,74,146,221,229,221,156,302,293,364,365,364,302,220,292,292,364,364,365,229,365,294,294,366,222,220,220,221,366,147,220,294,82,146,156,220,221,147,366,157,228,364,157,439,229,221,284,284,366,366,302,220,293,220,293,366,292,220,220,220,228,147,220,221,364,437,437,437,437,437,292,219,292,365,300,228,146,220,219,219,146,146,210,147,138,211,83,156,156,156,219,148,138,146,292,81,73,73,209,301,301,155,1,65,137,0,138,138,145,147,220,138,292,219,65,146,356,155,82,146,82,291,149,221,221,221,147,75,82,148,157,221,75,294,293,156,221,229,229,301,365,229,301,293,229,293,294,293,366,294,229,220,229,302,293,228,229,156,220,155,221,229,293,228,293,439,156,227,83,156,221,229,157,221,293,366,366,302,366,229,229,229,294,220,293,148,147,293,293,428,373,437,437,501,365,364,228,293,300,228,292,139,147,219,147,147,138,219,74,219,84,148,148,157,147,147,220,219,292,219,72,73,73,209,300,228,81,145,73,0,1,65,137,210,210,284,74,220,292,146,219,283,156,73,145,219,145,149,149,148,157,157,147,148,220,148,221,156,85,149,229,221,221,229,229,229,220,220,221,156,366,229,229,294,294,229,155,294,293,229,228,219,220,229,155,157,228,229,229,157,229,229,293,220,228,228,220,365,229,156,156,156,156,229,221,229,221,155,220,148,74,147,229,364,437,365,364,364,437,365,292,228,364,229,228,292,75,283,147,147,138,74,137,138,75,76,147,157,147,156,84,146,148,292,73,81,81,145,218,300,220,292,145,1,1,73,65,65,73,146,283,74,219,220,138,211,219,219,219,73,81,73,157,157,148,220,221,157,156,294,230,148,230,229,148,85,229,148,229,221,156,228,157,221,221,220,156,221,229,220,229,155,302,229,147,284,439,220,220,219,229,156,228,221,221,157,229,293,229,157,157,157,220,221,148,147,156,156,157,156,147,83,148,156,74,147,228,291,373,437,301,365,429,365,365,365,292,365,293,364,291,83,147,147,146,138,74,209,138,83,211,157,147,156,148,147,219,147,73,0,0,9,144,292,137,146,292,74,65,73,73,74,147,73,65,137,65,219,219,73,210,353,352,291,138,154,146,148,148,148,148,148,84,85,220,220,229,221,220,220,147,148,157,156,76,84,229,293,230,293,292,147,229,294,220,229,356,220,229,220,218,284,228,156,221,229,156,228,228,156,156,157,219,220,364,292,221,157,157,149,149,149,85,148,148,148,147,148,74,74,356,228,437,437,301,365,373,365,300,364,301,293,293,300,300,211,74,219,146,65,209,64,138,146,219,75,148,156,148,219,75,147,74,283,73,145,73,81,364,281,283,146,74,73,65,1,1,220,73,65,137,65,219,219,73,210,291,281,73,74,146,83,222,149,157,229,293,229,229,221,148,221,157,221,148,148,83,147,220,221,221,157,156,221,230,357,229,220,230,155,219,220,147,156,220,83,220,83,220,156,75,147,83,229,82,229,157,156,220,228,156,155,155,83,83,75,83,83,83,83,156,83,74,66,74,300,437,437,364,437,365,437,300,364,428,301,228,228,228,220,147,292,146,73,64,64,64,65,74,75,147,147,148,219,148,220,292,75,83,75,0,0,145,364,209,148,220,73,74,73,73,65,146,65,65,138,65,220,219,73,146,283,219,0,65,73,66,149,157,221,157,221,229,221,157,221,221,157,229,230,148,149,83,156,229,220,220,229,230,221,294,293,293,157,229,220,156,83,83,293,83,156,156,148,220,156,83,156,148,220,74,147,220,156,221,229,220,156,163,163,292,147,83,83,75,74,83,147,148,229,365,437,363,437,364,373,437,300,501,365,228,229,292,229,228,147,138,138,65,73,64,65,73,75,75,147,148,155,148,219,145,284,75,292,218,73,0,427,356,139,139,228,74,74,73,73,65,138,65,0,211,146,219,138,138,74,219,146,9,64,74,74,229,156,148,157,156,229,229,221,221,157,149,148,147,229,221,157,157,221,220,156,148,229,229,148,221,228,147,149,293,148,148,147,148,220,156,293,148,219,292,293,220,156,221,147,147,156,156,147,147,147,147,155,82,83,74,83,83,83,147,148,156,229,300,501,364,437,365,436,365,228,437,437,301,365,220,228,228,501,139,146,65,65,64,65,210,137,75,74,84,220,212,219,211,300,147,364,154,145,73,0,136,356,149,209,228,73,81,1,73,1,1,74,74,1,0,73,73,74,209,210,146,73,0,82,210,229,229,156,149,148,148,155,292,292,229,229,221,157,157,157,221,221,156,156,220,148,85,149,148,84,156,228,220,148,293,147,148,83,220,220,156,229,156,301,219,220,157,156,148,221,83,156,83,229,148,156,156,148,148,156,156,156,293,156,157,228,291,364,436,364,501,437,437,300,436,501,365,291,292,228,164,364,428,83,283,74,73,65,73,282,65,75,76,220,148,147,147,211,356,146,219,155,219,1,145,81,283,221,218,147,219,83,73,73,138,73,74,1,10,65,65,64,73,353,288,281,145,136,0,0,229,302,229,156,220,229,229,157,222,285,366,221,229,229,221,84,220,83,84,157,156,148,85,148,148,149,157,147,157,157,220,156,75,156,220,156,228,220,156,301,146,365,220,156,156,147,157,220,156,155,292,155,83,156,156,221,156,156,148,364,435,428,364,300,501,437,437,365,372,373,429,227,372,292,228,220,364,147,147,75,139,73,65,74,65,75,75,148,148,219,156,84,210,65,73,83,228,9,9,65,0,282,291,220,220,75,146,146,74,74,83,74,82,2,1,0,64,137,72,64,73,72,72,72,137,228,292,292,228,227,228,292,301,228,227,374,373,82,220,221,228,156,156,83,75,157,221,76,75,148,84,149,294,220,229,156,148,148,147,148,155,156,156,220,220,301,156,148,156,156,156,155,292,156,220,147,156,156,83,156,156,148,148,364,436,437,501,437,436,501,437,438,364,372,437,365,372,436,300,229,364,364,147,74,74,66,74,139,74,138,147,147,148,148,147,84,75,147,147,65,146,73,73,1,9,73,291,218,284,228,147,292,73,73,73,155,82,1,0,1,0,64,137,64,137,73,1,65,73,146,219,365,301,293,221,229,301,292,292,292,228,301,373,373,229,147,365,228,156,157,148,292,220,75,76,156,148,156,138,293,221,148,293,156,220,156,156,156,228,156,302,229,156,157,156,229,156,147,229,220,220,221,157,157,221,147,220,300,436,501,436,428,365,437,292,437,300,364,300,437,372,436,364,164,147,301,292,147,1,75,75,74,1,0,138,83,219,148,220,157,76,147,84,74,0,73,227,146,74,73,0,218,145,292,293,283,146,81,73,73,74,82,74,74,64,0,0,65,64,209,136,284,293,138,291,292,155,227

,300,293,301,301,301,301,229,301,373,364,228,219,229,229,300,301,228,156,148,147,156,148,76,83,156,148,147,301,148,84,156,220,229,301,220,220,156,220,301,228,157,293,229,157,156,147,156,83,156,157,220,156,228,437,437,437,227,292,437,501,437,228,428,373,228,501,365,364,364,228,156,228,301,292,74,138,138,65,1,137,65,147,211,148,147,221,76,147,84,74,147,138,65,218,74,0,73,9,283,209,364,292,219,81,1,66,1,74,146,74,73,74,74,64,64,136,201,136,284,221,73,291,228,292,300,364,364,364,427,364,364,364,364,373,373,373,300,292,220,229,292,374,364,292,220,82,292,221,292,148,157,148,138,293,148,156,156,157,221,229,293,292,221,366,301,157,157,220,229,157,221,148,83,229,220,221,229,365,428,429,228,437,437,437,364,437,501,364,300,437,364,436,292,228,228,147,301,292,219,138,74,1,65,65,64,73,146,148,84,147,84,147,76,75,148,83,219,146,73,81,82,81,73,356,217,355,291,73,66,2,64,137,145,73,74,74,1,0,65,0,137,201,136,293,293,1,291,300,372,300,300,364,364,301,373,373,437,436,436,364,155,220,301,219,147,156,220,228,364,220,221,228,300,220,74,220,292,157,229,220,149,156,156,156,156,229,292,156,221,220,229,221,156,156,229,229,220,147,156,147,221,228,428,228,437,501,501,501,429,437,437,509,428,428,437,436,228,228,228,219,219,300,227,291,282,0,0,1,64,64,74,147,148,148,148,147,148,147,156,76,211,147,210,74,220,74,9,73,136,217,209,219,210,67,74,137,146,73,74,74,0,0,0,137,137,137,200,137,292,293,65,283,364,363,372,300,373,364,437,437,437,437,437,436,381,363,364,227,373,155,147,156,220,292,292,229,221,228,364,156,83,284,157,156,229,220,157,156,156,156,221,156,220,157,156,302,221,156,221,221,302,221,220,364,220,229,227,437,437,501,501,355,437,428,501,509,364,437,437,437,292,300,364,436,147,301,291,436,218,64,65,65,137,64,64,65,75,76,219,76,220,147,148,76,83,147,74,73,292,74,81,81,73,218,138,75,74,73,138,292,82,147,146,73,1,74,74,73,72,65,137,201,146,292,292,65,283,299,372,372,436,436,435,436,435,435,363,436,373,381,435,508,436,227,373,364,301,147,147,292,156,148,221,227,365,221,149,149,84,156,147,156,221,156,221,220,156,220,220,157,301,229,429,220,229,301,221,356,220,229,228,437,437,501,437,364,501,437,501,437,501,501,437,437,437,373,364,436,219,292,365,301,364,73,74,210,64,73,0,73,0,76,76,3,148,76,75,76,76,147,74,210,146,147,81,292,81,291,283,75,355,74,75,82,74,147,210,83,83,74,136,0,0,0,137,137,137,146,292,356,64,283,436,436,436,372,436,508,499,499,507,499,499,499,362,437,437,436,435,155,156,147,300,219,156,156,221,148,229,218,292,157,221,157,156,156,229,229,221,221,221,155,147,228,156,301,157,293,229,229,220,156,156,228,365,437,364,437,364,292,437,437,437,437,436,437,373,437,437,364,372,436,292,82,372,292,292,501,0,138,74,1,65,65,74,0,75,75,76,76,147,147,84,75,220,146,138,365,73,228,73,73,81,75,218,74,75,81,146,74,219,147,210,74,73,0,10,2,0,73,137,136,137,356,219,0,209,436,364,436,444,435,435,499,435,499,508,508,427,435,228,218,372,300,435,156,156,229,300,155,74,147,157,148,220,292,229,221,10,148,147,148,229,156,220,156,293,156,228,221,229,229,293,229,156,221,156,229,365,437,437,437,428,365,365,437,437,364,437,437,373,428,437,364,372,364,292,147,364,228,228,364,427,0,66,74,1,0,65,1,0,138,76,75,83,147,84,75,147,147,201,1,146,292,73,218,73,73,147,211,75,74,75,146,74,146,155,137,74,1,74,137,0,65,137,73,0,1,65,65,73,73,436,363,436,435,435,435,499,435,444,435,427,435,499,508,436,228,436,373,436,228,156,292,155,219,146,365,221,221,293,220,221,229,148,147,220,148,302,148,220,156,229,221,221,229,221,229,229,221,148,293,365,437,437,437,437,292,301,372,300,364,429,373,373,437,437,292,372,436,292,220,219,363,220,82,428,137,65,75,1,0,65,1,138,0,75,75,84,148,148,75,147,147,75,75,65,74,82,146,148,283,73,283,75,74,76,218,73,73,211,147,82,146,74,138,74,74,138,64,137,209,0,209,73,210,292,372,435,508,436,437,501,509,427,500,500,500,436,434,435,500,444,373,436,436,436,156,147,373,219,291,373,292,220,291,156,292,157,148,147,292,221,229,156,148,148,365,156,221,229,220,293,156,156,157,429,428,501,435,364,437,365,437,228,365,428,372,228,428,365,437,437,291,292,220,219,364,300,220,364,364,65,65,65,138,1,65,74,73,65,220,76,219,147,147,147,147,75,147,74,1,65,300,74,82,74,137,290,146,75,74,217,138,74,73,147,228,146,66,228,82,65,74,1,65,1,0,72,137,219,284,435,435,500,500,500,508,508,508,436,500,500,500,435,508,435,436,372,436,372,437,427,291,364,373,219,429,364,292,221,220,229,221,156,156,293,293,156,229,148,157,301,148,220,229,157,220,156,156,365,356,429,436,364,437,373,428,365,429,501,227,228,364,365,437,437,437,228,219,283,428,365,300,292,364,219,0,1,74,65,66,65,65,64,219,76,148,148,84,147,147,75,147,147,75,146,0,73,82,64,82,209,209,137,210,138,291,83,81,137,137,219,65,163,219,66,219,74,1,9,10,0,8,0,211,219,436,435,435,499,434,426,427,435,435,499,435,508,508,435,435,435,436,362,435,363,436,364,427,372,437,283,362,156,148,219,221,156,221,157,220,293,220,156,229,157,229,147,221,229,156,221,221,156,365,364,501,436,429,437,365,437,437,501,364,228,292,437,501,437,291,292,228,291,364,292,292,364,228,228,219,74,66,65,65,1,0,0,146,76,147,220,76,147,147,66,219,139,147,211,218,82,283,81,74,73,139,209,72,218,147,147,137,145,73,291,146,82,228,219,219,146,73,137,137,137,0,72,0,64,0,436,499,499,435,490,489,489,424,489,353,426,500,508,499,500,435,499,436,363,435,434,436,292,434,501,300,428,293,156,156,220,156,221,157,84,221,221,148,147,221,220,229,220,220,156,220,220,293,364,428,427,429,501,435,501,501,436,292,228,300,363,437,429,228,228,292,364,220,228,228,364,220,228,364,218,73,0,1,65,66,0,65,76,147,212,76,147,147,155,156,147,147,220,219,73,292,72,0,73,72,75,210,137,138,91,75,137,74,83,74,74,218,145,292,219,147,73,1,0,0,0,73,64,210,0,508,435,435,489,489,489,497,489,489,489,416,489,435,508,427,508,426,508,435,436,426,426,437,364,499,364,155,354,83,221,155,293,157,293,84,148,230,148,156,229,229,221,156,156,220,229,221,365,356,427,500,437,435,501,501,436,291,364,365,364,501,283,293,228,365,436,155,292,220,228,228,220,292,364,145,0,1,2,65,73,65,147,147,147,148,75,148,147,147,147,147,155,156,219,291,145,218,72,73,291,147,209,138,83,146,146,155,73,73,82,83,82,73,138,291,145,9,82,138,73,64,81,64,146,74,435,425,489,497,489,489,489,489,489,489,489,416,489,435,499,435,508,426,499,435,373,354,436,373,292,428,364,364,220,221,292,157,221,221,156,157,220,148,220,293,229,229,221,156,221,293,229,366,365,363,365,363,364,501,428,428,365,364,437,365,291,292,364,437,363,156,292,219,291,292,228,364,428,428,0,1,1,74,65,65,138,147,220,147,83,148,84,76,156,220,155,75,220,292,365,301,292,81,218,363,146,145,74,138,73,219,73,73,83,74,1,73,73,73,300,147,147,73,65,73,64,64,65,146,283,489,497,489,489,489,489,489,489,489,489,489,489,489,489,425,435,499,498,435,499,436,437,426,437,437,291,292,283,148,156,228,148,221,221,220,157,221,148,156,229,221,229,221,220,221,156,293,302,365,429,301,435,501,501,354,365,365,364,364,291,228,364,364,292,147,220,364,147,292,364,72,65,0,0,0,74,2,2,73,65,84,147,147,147,147,147,148,147,76,220,75,220,147,76,219,373,73,148,147,282,291,145,147,138,292,292,219,220,73,73,218,73,73,72,228,73,147,10,0,137,0,0,65,146,219,489,425,489,489,489,488,489,489,489,497,489,425,489,489,489,416,435,508,500,353,499,435,500,434,373,300,228,155,156,148,221,229,157,229,292,221,221,148,147,229,148,229,157,220,220,220,302,366,429,366,428,428,437,362,301,365,429,437,364,292,364,365,292,219,156,364,156,292,364,72,0,0,65,0,1,2,65,73,73,146,148,148,84,147,147,219,155,76,293,148,293,76,220,211,227,73,82,218,82,82,290,209,146,210,300,154,228,219,146,227,74,73,146,137,219,138,74,0,0,0,0,65,0,146,219,425,489,489,489,489,489,489,489,489,489,425,416,489,425,425,489,345,436,499,508,426,435,292,490,437,373,156,300,228,221,148,301,157,156,148,147,156,147,83,221,147,229,220,220,293,229,302,365,365,365,365,429,435,363,365,365,429,429,364,365,364,155,83,220,292,155,228,364,492,0,0,75,74,74,0,73,1,1,0,148,155,76,155,219,147,147,148,220,220,148,220,220,284,75,210,65,219,146,81,81,210,218,282,282,292,219,220,146,291,219,218,73,138,65,138,65,1,0,0,0,219,138,137,211,219,425,489,425,425,417,489,424,489,489,489,489,489,425,425,416,416,425,363,500,435,353,499,364,364,499,373,373,220,164,157,221,300,221,221,148,156,156,220,148,221,155,156,156,147,293,229,366,366,437,365,365,428,434,365,365,437,364,364,365,365,365,219,292,220,147,292,156,219,218,0,75,74,66,65,65,65,65,138,65,291,76,147,219,147,147,220,220,219,148,220,220,220,75,219,282,219,73,147,75,146,145,291,291,210,137,228,228,146,147,146,146,74,219,1,1,0,0,0,73,65,211,74,137,210,211,489,417

,426,499,499,499,499,489,489,489,489,425,489,425,416,416,416,417,426,435,362,435,364,437,437,372,300,229,164,221,219,219,221,221,156,156,221,148,84,221,148,148,156,83,220,293,293,437,364,365,437,427,428,365,364,437,501,437,365,364,365,300,292,156,292,219,155,219,64,0,74,74,65,64,0,73,1,65,138,219,148,220,148,84,147,219,147,75,148,219,148,147,220,75,138,137,65,145,81,81,209,282,355,211,66,219,219,219,219,218,146,146,138,0,1,1,0,0,65,65,219,66,64,137,0,416,499,500,499,499,499,499,499,499,490,489,425,425,425,416,425,425,416,426,499,435,435,435,427,437,364,364,301,228,229,147,155,156,156,156,155,221,147,84,228,156,156,220,156,157,293,365,501,365,437,428,363,437,365,437,429,501,365,365,365,365,156,292,364,219,228,155,147,73,0,64,66,65,65,65,1,74,73,210,148,156,147,75,219,147,148,147,147,147,220,211,156,75,75,291,81,73,64,73,73,145,218,355,66,74,137,211,138,147,146,146,292,146,1,64,65,0,1,65,137,211,75,65,73,72,499,500,499,498,499,499,435,499,435,499,498,489,425,497,489,416,425,425,418,499,435,435,435,500,500,364,364,364,228,365,157,156,147,156,147,220,157,220,148,228,220,157,219,221,229,428,429,364,428,437,427,437,501,427,437,501,429,365,429,365,220,292,364,219,219,355,147,219,64,0,74,65,65,1,74,73,65,65,210,220,219,76,147,147,76,83,147,147,292,219,148,148,220,292,147,81,81,145,145,81,209,283,282,66,73,66,145,73,74,219,146,146,64,356,137,0,0,65,65,219,146,75,137,65,81,500,434,435,499,499,500,499,499,427,426,499,498,489,416,425,425,425,425,344,435,435,435,499,363,436,509,427,363,292,365,229,157,156,155,220,155,220,156,221,220,156,156,155,229,292,364,428,501,436,428,500,501,436,364,428,501,437,501,364,292,228,364,300,292,218,227,219,219,0,0,1,66,65,65,1,1,1,64,211,219,148,155,219,84,147,147,219,220,147,156,220,292,220,75,220,219,283,137,64,217,146,291,145,74,209,138,81,147,146,74,146,145,73,291,73,65,0,0,65,210,137,75,65,219,81,499,499,427,435,436,435,435,436,435,426,426,499,489,425,425,425,490,416,417,499,435,435,435,363,364,436,355,147,218,292,156,148,156,292,220,156,292,156,221,156,147,156,156,291,291,428,500,437,428,501,501,363,428,437,437,364,501,437,364,292,364,292,428,73,65,218,219,427,0,64,65,1,1,0,0,0,0,0,211,219,220,219,83,83,146,219,147,220,147,293,292,212,76,220,211,292,145,208,144,209,74,291,145,219,210,138,73,219,146,74,81,73,0,146,74,1,0,0,0,211,138,75,73,291,65,435,500,435,426,426,426,427,361,435,435,499,435,490,425,417,417,425,425,425,500,435,500,434,300,373,363,219,83,219,292,156,84,156,211,156,155,292,156,220,220,148,156,156,219,219,427,501,428,501,501,364,363,437,437,364,501,436,437,291,364,364,364,363,65,64,64,363,210,0,0,0,64,0,0,0,0,0,65,138,147,211,219,147,213,211,147,210,219,219,284,76,76,220,76,284,137,217,216,144,209,75,282,209,283,145,219,146,82,73,82,73,81,0,73,9,0,1,64,0,146,147,65,292,219,136,435,435,435,435,426,434,426,499,426,435,500,435,499,425,489,425,417,344,428,500,499,499,435,291,364,437,363,83,365,228,155,147,156,147,147,156,156,156,284,147,148,156,148,292,219,428,364,436,436,435,364,437,437,364,437,501,429,429,429,292,364,219,428,0,0,0,1,1,0,0,0,0,65,0,0,64,73,0,291,75,219,147,147,211,147,147,211,219,219,75,146,220,84,75,146,72,216,74,209,145,145,291,282,291,218,291,146,64,1,1,73,73,137,73,209,65,65,0,0,219,146,65,291,137,137,500,435,499,435,435,500,499,499,426,499,426,435,490,425,425,489,344,344,436,508,499,500,499,291,364,365,363,220,300,220,220,148,156,147,147,155,155,147,220,74,148,156,148,219,291,364,428,501,427,363,364,437,364,428,501,364,437,428,292,292,292,156,428,0,136,0,0,0,64,0,0,1,0,73,64,0,0,0,220,83,147,76,147,147,76,147,147,219,147,219,220,76,147,147,139,64,208,74,218,218,144,217,291,363,283,0,65,0,0,0,0,64,292,73,137,65,1,0,65,211,210,0,219,201,73,435,435,434,435,426,426,499,435,435,499,498,426,425,417,425,489,416,344,435,500,500,436,427,300,292,291,292,292,220,229,147,147,156,220,147,220,155,138,155,138,156,229,156,219,364,364,364,364,427,428,501,364,428,501,291,437,437,220,220,364,156,356,218,72,64,0,0,0,0,0,0,1,64,65,1,65,65,0,75,219,219,147,219,76,147,75,219,76,219,148,148,219,148,76,420,64,73,210,283,210,283,145,290,209,137,1,138,81,81,9,0,1,218,73,137,0,65,73,65,211,210,64,65,73,73,436,435,426,426,427,427,426,498,435,435,435,426,426,425,417,490,490,416,499,299,436,435,364,435,363,218,301,228,147,220,155,73,83,228,147,220,220,74,147,74,156,229,220,283,363,428,427,427,437,501,363,428,437,437,437,437,292,228,364,292,292,492,64,0,64,0,0,0,0,0,0,64,64,0,0,0,65,64,292,147,147,211,76,148,76,147,76,211,147,138,147,212,75,219,148,72,137,217,219,64,282,137,218,137,1,73,73,9,73,9,73,146,73,83,73,65,1,0,138,64,209,284,64,137,137,426,427,362,427,435,435,434,435,434,427,426,426,426,425,489,417,408,435,435,363,436,364,364,373,229,226,364,221,156,147,83,73,83,220,228,221,219,283,147,74,156,156,292,428,363,363,436,428,428,363,427,437,437,437,437,364,292,364,429,292,428,427,65,64,0,0,0,0,0,0,0,1,65,0,1,1,1,65,219,75,147,75,75,147,147,147,211,147,148,75,219,147,147,75,137,0,72,144,218,73,283,145,218,73,74,146,1,227,73,1,1,218,73,83,81,65,0,64,73,138,146,283,65,64,65,427,427,362,363,363,363,427,427,435,426,425,361,416,425,416,344,416,363,364,364,508,226,373,373,220,292,227,157,148,220,292,73,156,291,156,155,221,155,138,73,156,220,356,363,362,364,364,437,355,363,501,437,437,428,437,292,364,364,291,428,428,146,145,64,0,0,0,0,0,64,1,65,0,1,0,0,137,64,219,147,147,147,219,146,219,147,147,76,75,219,147,146,147,138,1,218,136,137,209,146,209,218,209,146,364,73,291,81,9,146,73,145,74,83,73,0,0,73,65,146,146,147,65,65,0,427,354,427,426,362,290,362,427,427,362,426,408,416,416,408,416,435,436,363,436,436,300,437,364,292,365,164,156,156,157,155,147,221,219,157,220,221,146,74,147,156,220,290,363,363,435,355,283,292,501,428,437,428,428,292,364,364,228,364,429,428,73,0,0,0,0,1,137,0,0,1,1,0,65,1,1,73,73,75,211,147,147,74,147,219,147,147,138,146,147,74,147,147,65,73,72,145,72,209,209,218,145,64,73,219,0,219,73,283,147,74,74,74,83,9,0,0,0,73,146,210,211,74,65,1,364,427,427,219,364,363,362,435,354,426,353,344,408,417,427,436,364,435,436,364,299,300,427,219,427,291,365,220,156,156,220,147,147,228,156,83,156,146,73,147,219,292,435,363,437,291,292,355,437,364,437,428,436,355,292,364,228,228,364,428,218,64,0,0,0,64,65,0,64,0,0,0,65,65,0,0,65,64,219,75,147,74,74,219,147,147,146,83,147,146,147,147,146,73,145,218,138,210,218,72,282,65,73,64,65,219,219,0,218,65,146,138,74,82,9,73,1,0,65,74,210,139,1,0,65,300,291,363,435,436,435,363,363,417,417,417,363,372,364,373,299,435,363,436,301,299,364,364,292,146,292,220,156,155,147,220,219,147,228,74,147,155,147,83,147,228,364,363,437,428,364,428,501,291,364,428,364,364,356,364,291,292,364,364,356,146,64,0,0,0,0,0,65,73,0,0,0,0,0,0,0,65,73,211,147,146,74,147,147,83,146,76,147,147,147,147,146,146,137,137,218,73,283,218,73,218,137,210,72,72,218,291,73,219,73,82,146,65,82,73,0,1,0,64,146,210,75,1,0,147,300,300,291,363,363,435,436,436,291,299,363,363,435,373,219,435,364,221,301,363,435,373,227,219,146,219,83,227,146,156,156,156,220,220,147,147,227,221,147,147,220,363,436,428,363,428,292,428,429,364,364,356,292,219,428,292,365,364,228,364,73,0,0,0,64,65,1,1,65,65,0,0,0,1,66,65,146,73,211,138,74,147,147,83,146,147,147,147,147,147,146,147,146,73,65,282,137,136,217,73,209,218,138,66,0,72,0,146,210,73,219,355,73,74,74,0,1,0,1,64,209,66,0,147,147,428,291,362,427,291,219,227,227,363,363,291,363,364,301,364,364,437,219,291,435,372,227,219,292,220,219,83,155,155,156,156,156,164,219,156,156,147,146,147,219,292,363,437,363,428,364,364,428,292,364,364,292,219,364,291,291,364,220,292,428,74,0,0,65,0,0,0,1,137,0,0,0,1,65,65,1,138,0,219,74,147,211,74,147,146,146,147,84,147,147,75,74,75,74,65,210,145,72,218,137,72,282,74,219,1,1,1,145,146,74,292,74,73,210,73,65,0,0,0,0,209,74,1,74,74,220,355,363,427,362,427,427,364,364,364,364,363,309,300,364,372,291,228,427,364,146,228,300,292,155,219,156,219,155,147,156,155,228,73,156,83,156,138,147,219,363,436,355,364,363,292,437,365,364,428,292,364,364,364,428,364,300,155,292,364,146,73,0,0,0,0,65,64,65,1,65,1,0,0,0,0,65,0,146,10,219,74,147,146,74,74,146,146,146,75,75,147,75,74,138,72,145,144,137,145,210,72,74,210,0,137,0,0,0,74,292,73,73,146,73,0,0,0,1,73,137,66,0,74,147,291,300,300,300,365,299,227,291,363,427,363,300,291,300,300,227,364,300,436,291,147,220,300,156,147,156,156,155,219,219,155,155,219,82,220,155,147,82,362,219,428,428,364,436,292,437,364,356,428,291,356,219,364,355,364,364,220,428,228,364,291,0,0,0,0,73,0,74,74,65,0,0,0,0,0,0,1,1,66,74,147,74,211,74,66,74,146,146,75,75,138,76,146,65,73,73,209,136,209,137,209,145,210,282,72,64,0,0,0,138,146,146,73,146,65,65,0,1,0,0,0,66,1,74,147};
		logic [23:0] idx;
		assign idx = (nX/2)*125 + (nY/2);
		assign cidx = IMG[24999 - idx];
		
endmodule
